module sbtm_a0 (input  logic [6:0] a,
		output logic [12:0] y);
   always_comb
     case(a)
       7'b0000000: y = 13'b1111111100010;
       7'b0000001: y = 13'b1111110100011;
       7'b0000010: y = 13'b1111101100101;
       7'b0000011: y = 13'b1111100101000;
       7'b0000100: y = 13'b1111011101100;
       7'b0000101: y = 13'b1111010110000;
       7'b0000110: y = 13'b1111001110110;
       7'b0000111: y = 13'b1111000111100;
       7'b0001000: y = 13'b1111000000100;
       7'b0001001: y = 13'b1110111001100;
       7'b0001010: y = 13'b1110110010101;
       7'b0001011: y = 13'b1110101011110;
       7'b0001100: y = 13'b1110100101001;
       7'b0001101: y = 13'b1110011110100;
       7'b0001110: y = 13'b1110011000000;
       7'b0001111: y = 13'b1110010001101;
       7'b0010000: y = 13'b1110001011010;
       7'b0010001: y = 13'b1110000101000;
       7'b0010010: y = 13'b1101111110111;
       7'b0010011: y = 13'b1101111000110;
       7'b0010100: y = 13'b1101110010111;
       7'b0010101: y = 13'b1101101100111;
       7'b0010110: y = 13'b1101100111001;
       7'b0010111: y = 13'b1101100001011;
       7'b0011000: y = 13'b1101011011101;
       7'b0011001: y = 13'b1101010110001;
       7'b0011010: y = 13'b1101010000100;
       7'b0011011: y = 13'b1101001011001;
       7'b0011100: y = 13'b1101000101110;
       7'b0011101: y = 13'b1101000000011;
       7'b0011110: y = 13'b1100111011001;
       7'b0011111: y = 13'b1100110101111;
       7'b0100000: y = 13'b1100110000110;
       7'b0100001: y = 13'b1100101011110;
       7'b0100010: y = 13'b1100100110110;
       7'b0100011: y = 13'b1100100001111;
       7'b0100100: y = 13'b1100011101000;
       7'b0100101: y = 13'b1100011000001;
       7'b0100110: y = 13'b1100010011011;
       7'b0100111: y = 13'b1100001110101;
       7'b0101000: y = 13'b1100001010000;
       7'b0101001: y = 13'b1100000101011;
       7'b0101010: y = 13'b1100000000111;
       7'b0101011: y = 13'b1011111100011;
       7'b0101100: y = 13'b1011111000000;
       7'b0101101: y = 13'b1011110011101;
       7'b0101110: y = 13'b1011101111010;
       7'b0101111: y = 13'b1011101011000;
       7'b0110000: y = 13'b1011100110110;
       7'b0110001: y = 13'b1011100010101;
       7'b0110010: y = 13'b1011011110011;
       7'b0110011: y = 13'b1011011010011;
       7'b0110100: y = 13'b1011010110010;
       7'b0110101: y = 13'b1011010010010;
       7'b0110110: y = 13'b1011001110011;
       7'b0110111: y = 13'b1011001010011;
       7'b0111000: y = 13'b1011000110100;
       7'b0111001: y = 13'b1011000010110;
       7'b0111010: y = 13'b1010111110111;
       7'b0111011: y = 13'b1010111011001;
       7'b0111100: y = 13'b1010110111100;
       7'b0111101: y = 13'b1010110011110;
       7'b0111110: y = 13'b1010110000001;
       7'b0111111: y = 13'b1010101100100;
       7'b1000000: y = 13'b1010101001000;
       7'b1000001: y = 13'b1010100101100;
       7'b1000010: y = 13'b1010100010000;
       7'b1000011: y = 13'b1010011110100;
       7'b1000100: y = 13'b1010011011001;
       7'b1000101: y = 13'b1010010111110;
       7'b1000110: y = 13'b1010010100011;
       7'b1000111: y = 13'b1010010001001;
       7'b1001000: y = 13'b1010001101111;
       7'b1001001: y = 13'b1010001010101;
       7'b1001010: y = 13'b1010000111011;
       7'b1001011: y = 13'b1010000100001;
       7'b1001100: y = 13'b1010000001000;
       7'b1001101: y = 13'b1001111101111;
       7'b1001110: y = 13'b1001111010111;
       7'b1001111: y = 13'b1001110111110;
       7'b1010000: y = 13'b1001110100110;
       7'b1010001: y = 13'b1001110001110;
       7'b1010010: y = 13'b1001101110110;
       7'b1010011: y = 13'b1001101011111;
       7'b1010100: y = 13'b1001101000111;
       7'b1010101: y = 13'b1001100110000;
       7'b1010110: y = 13'b1001100011001;
       7'b1010111: y = 13'b1001100000010;
       7'b1011000: y = 13'b1001011101100;
       7'b1011001: y = 13'b1001011010110;
       7'b1011010: y = 13'b1001011000000;
       7'b1011011: y = 13'b1001010101010;
       7'b1011100: y = 13'b1001010010100;
       7'b1011101: y = 13'b1001001111111;
       7'b1011110: y = 13'b1001001101001;
       7'b1011111: y = 13'b1001001010100;
       7'b1100000: y = 13'b1001000111111;
       7'b1100001: y = 13'b1001000101011;
       7'b1100010: y = 13'b1001000010110;
       7'b1100011: y = 13'b1001000000010;
       7'b1100100: y = 13'b1000111101110;
       7'b1100101: y = 13'b1000111011010;
       7'b1100110: y = 13'b1000111000110;
       7'b1100111: y = 13'b1000110110010;
       7'b1101000: y = 13'b1000110011111;
       7'b1101001: y = 13'b1000110001011;
       7'b1101010: y = 13'b1000101111000;
       7'b1101011: y = 13'b1000101100101;
       7'b1101100: y = 13'b1000101010010;
       7'b1101101: y = 13'b1000101000000;
       7'b1101110: y = 13'b1000100101101;
       7'b1101111: y = 13'b1000100011011;
       7'b1110000: y = 13'b1000100001001;
       7'b1110001: y = 13'b1000011110110;
       7'b1110010: y = 13'b1000011100101;
       7'b1110011: y = 13'b1000011010011;
       7'b1110100: y = 13'b1000011000001;
       7'b1110101: y = 13'b1000010110000;
       7'b1110110: y = 13'b1000010011110;
       7'b1110111: y = 13'b1000010001101;
       7'b1111000: y = 13'b1000001111100;
       7'b1111001: y = 13'b1000001101011;
       7'b1111010: y = 13'b1000001011010;
       7'b1111011: y = 13'b1000001001010;
       7'b1111100: y = 13'b1000000111001;
       7'b1111101: y = 13'b1000000101001;
       7'b1111110: y = 13'b1000000011001;
       7'b1111111: y = 13'b1000000001001;	    
       default: y = 13'bxxxxxxxxxxxxx;
     endcase // case (a)
    
endmodule // sbtm_a0
// This module implements a 52-bit carry lookahead adder. It is used
// for rounding in the floating point adder. 

module cla52 (S, CO, X, Y);
   
   input  [51:0] X;
   input [51:0]  Y;
   
   output [51:0] S;
   output 	 CO;
   
   wire [63:0] 	 A,B,Q;//***KEP was 0:63 - changed due to lint warning
   wire 	 LOGIC0;
   wire 	 CIN;
   wire 	 CO_64;
   
   assign LOGIC0 = 0;
   assign CIN = 0;
   DBLCADDER_64_64 U1 (A , B , CIN, Q , CO_64);
   assign A[0] = X[0];
   assign B[0] = Y[0];
   assign A[1] = X[1];
   assign B[1] = Y[1];
   assign A[2] = X[2];
   assign B[2] = Y[2];
   assign A[3] = X[3];
   assign B[3] = Y[3];
   assign A[4] = X[4];
   assign B[4] = Y[4];
   assign A[5] = X[5];
   assign B[5] = Y[5];
   assign A[6] = X[6];
   assign B[6] = Y[6];
   assign A[7] = X[7];
   assign B[7] = Y[7];
   assign A[8] = X[8];
   assign B[8] = Y[8];
   assign A[9] = X[9];
   assign B[9] = Y[9];
   assign A[10] = X[10];
   assign B[10] = Y[10];
   assign A[11] = X[11];
   assign B[11] = Y[11];
   assign A[12] = X[12];
   assign B[12] = Y[12];
   assign A[13] = X[13];
   assign B[13] = Y[13];
   assign A[14] = X[14];
   assign B[14] = Y[14];
   assign A[15] = X[15];
   assign B[15] = Y[15];
   assign A[16] = X[16];
   assign B[16] = Y[16];
   assign A[17] = X[17];
   assign B[17] = Y[17];
   assign A[18] = X[18];
   assign B[18] = Y[18];
   assign A[19] = X[19];
   assign B[19] = Y[19];
   assign A[20] = X[20];
   assign B[20] = Y[20];
   assign A[21] = X[21];
   assign B[21] = Y[21];
   assign A[22] = X[22];
   assign B[22] = Y[22];
   assign A[23] = X[23];
   assign B[23] = Y[23];
   assign A[24] = X[24];
   assign B[24] = Y[24];
   assign A[25] = X[25];
   assign B[25] = Y[25];
   assign A[26] = X[26];
   assign B[26] = Y[26];
   assign A[27] = X[27];
   assign B[27] = Y[27];
   assign A[28] = X[28];
   assign B[28] = Y[28];
   assign A[29] = X[29];
   assign B[29] = Y[29];
   assign A[30] = X[30];
   assign B[30] = Y[30];
   assign A[31] = X[31];
   assign B[31] = Y[31];
   assign A[32] = X[32];
   assign B[32] = Y[32];
   assign A[33] = X[33];
   assign B[33] = Y[33];
   assign A[34] = X[34];
   assign B[34] = Y[34];
   assign A[35] = X[35];
   assign B[35] = Y[35];
   assign A[36] = X[36];
   assign B[36] = Y[36];
   assign A[37] = X[37];
   assign B[37] = Y[37];
   assign A[38] = X[38];
   assign B[38] = Y[38];
   assign A[39] = X[39];
   assign B[39] = Y[39];
   assign A[40] = X[40];
   assign B[40] = Y[40];
   assign A[41] = X[41];
   assign B[41] = Y[41];
   assign A[42] = X[42];
   assign B[42] = Y[42];
   assign A[43] = X[43];
   assign B[43] = Y[43];
   assign A[44] = X[44];
   assign B[44] = Y[44];
   assign A[45] = X[45];
   assign B[45] = Y[45];
   assign A[46] = X[46];
   assign B[46] = Y[46];
   assign A[47] = X[47];
   assign B[47] = Y[47];
   assign A[48] = X[48];
   assign B[48] = Y[48];
   assign A[49] = X[49];
   assign B[49] = Y[49];
   assign A[50] = X[50];
   assign B[50] = Y[50];
   assign A[51] = X[51];
   assign B[51] = Y[51];
   assign A[52] = LOGIC0;
   assign B[52] = LOGIC0;
   assign A[53] = LOGIC0;
   assign B[53] = LOGIC0;
   assign A[54] = LOGIC0;
   assign B[54] = LOGIC0;
   assign A[55] = LOGIC0;
   assign B[55] = LOGIC0;
   assign A[56] = LOGIC0;
   assign B[56] = LOGIC0;
   assign A[57] = LOGIC0;
   assign B[57] = LOGIC0;
   assign A[58] = LOGIC0;
   assign B[58] = LOGIC0;
   assign A[59] = LOGIC0;
   assign B[59] = LOGIC0;
   assign A[60] = LOGIC0;
   assign B[60] = LOGIC0;
   assign A[61] = LOGIC0;
   assign B[61] = LOGIC0;
   assign A[62] = LOGIC0;
   assign B[62] = LOGIC0;
   assign A[63] = LOGIC0;
   assign B[63] = LOGIC0;
   assign S[0] = Q[0];
   assign S[1] = Q[1];
   assign S[2] = Q[2];
   assign S[3] = Q[3];
   assign S[4] = Q[4];
   assign S[5] = Q[5];
   assign S[6] = Q[6];
   assign S[7] = Q[7];
   assign S[8] = Q[8];
   assign S[9] = Q[9];
   assign S[10] = Q[10];
   assign S[11] = Q[11];
   assign S[12] = Q[12];
   assign S[13] = Q[13];
   assign S[14] = Q[14];
   assign S[15] = Q[15];
   assign S[16] = Q[16];
   assign S[17] = Q[17];
   assign S[18] = Q[18];
   assign S[19] = Q[19];
   assign S[20] = Q[20];
   assign S[21] = Q[21];
   assign S[22] = Q[22];
   assign S[23] = Q[23];
   assign S[24] = Q[24];
   assign S[25] = Q[25];
   assign S[26] = Q[26];
   assign S[27] = Q[27];
   assign S[28] = Q[28];
   assign S[29] = Q[29];
   assign S[30] = Q[30];
   assign S[31] = Q[31];
   assign S[32] = Q[32];
   assign S[33] = Q[33];
   assign S[34] = Q[34];
   assign S[35] = Q[35];
   assign S[36] = Q[36];
   assign S[37] = Q[37];
   assign S[38] = Q[38];
   assign S[39] = Q[39];
   assign S[40] = Q[40];
   assign S[41] = Q[41];
   assign S[42] = Q[42];
   assign S[43] = Q[43];
   assign S[44] = Q[44];
   assign S[45] = Q[45];
   assign S[46] = Q[46];
   assign S[47] = Q[47];
   assign S[48] = Q[48];
   assign S[49] = Q[49];
   assign S[50] = Q[50];
   assign S[51] = Q[51];
   assign CO    = Q[52];
   
endmodule //cla52

// This module implements a 52-bit carry lookahead subtractor. It is used
// for rounding in the floating point adder. 

module cla_sub52 (S, X, Y);
   
   input [51:0] X;
   input [51:0] Y;
   
   output [51:0] S;
   
   wire [63:0] 	 A,B,Q,Bbar;//***KEP was 0:63 - changed due to lint warning
   wire 	 LOGIC0;
   wire 	 CIN;
   wire 	 CO_52;
   wire   CO_64;
   
   assign Bbar = ~B;
   assign LOGIC0 = 0;
   assign CIN = 0;

   DBLCADDER_64_64 U1 (A , Bbar , CIN, Q , CO_64);

   assign A[0] = X[0];
   assign B[0] = Y[0];
   assign A[1] = X[1];
   assign B[1] = Y[1];
   assign A[2] = X[2];
   assign B[2] = Y[2];
   assign A[3] = X[3];
   assign B[3] = Y[3];
   assign A[4] = X[4];
   assign B[4] = Y[4];
   assign A[5] = X[5];
   assign B[5] = Y[5];
   assign A[6] = X[6];
   assign B[6] = Y[6];
   assign A[7] = X[7];
   assign B[7] = Y[7];
   assign A[8] = X[8];
   assign B[8] = Y[8];
   assign A[9] = X[9];
   assign B[9] = Y[9];
   assign A[10] = X[10];
   assign B[10] = Y[10];
   assign A[11] = X[11];
   assign B[11] = Y[11];
   assign A[12] = X[12];
   assign B[12] = Y[12];
   assign A[13] = X[13];
   assign B[13] = Y[13];
   assign A[14] = X[14];
   assign B[14] = Y[14];
   assign A[15] = X[15];
   assign B[15] = Y[15];
   assign A[16] = X[16];
   assign B[16] = Y[16];
   assign A[17] = X[17];
   assign B[17] = Y[17];
   assign A[18] = X[18];
   assign B[18] = Y[18];
   assign A[19] = X[19];
   assign B[19] = Y[19];
   assign A[20] = X[20];
   assign B[20] = Y[20];
   assign A[21] = X[21];
   assign B[21] = Y[21];
   assign A[22] = X[22];
   assign B[22] = Y[22];
   assign A[23] = X[23];
   assign B[23] = Y[23];
   assign A[24] = X[24];
   assign B[24] = Y[24];
   assign A[25] = X[25];
   assign B[25] = Y[25];
   assign A[26] = X[26];
   assign B[26] = Y[26];
   assign A[27] = X[27];
   assign B[27] = Y[27];
   assign A[28] = X[28];
   assign B[28] = Y[28];
   assign A[29] = X[29];
   assign B[29] = Y[29];
   assign A[30] = X[30];
   assign B[30] = Y[30];
   assign A[31] = X[31];
   assign B[31] = Y[31];
   assign A[32] = X[32];
   assign B[32] = Y[32];
   assign A[33] = X[33];
   assign B[33] = Y[33];
   assign A[34] = X[34];
   assign B[34] = Y[34];
   assign A[35] = X[35];
   assign B[35] = Y[35];
   assign A[36] = X[36];
   assign B[36] = Y[36];
   assign A[37] = X[37];
   assign B[37] = Y[37];
   assign A[38] = X[38];
   assign B[38] = Y[38];
   assign A[39] = X[39];
   assign B[39] = Y[39];
   assign A[40] = X[40];
   assign B[40] = Y[40];
   assign A[41] = X[41];
   assign B[41] = Y[41];
   assign A[42] = X[42];
   assign B[42] = Y[42];
   assign A[43] = X[43];
   assign B[43] = Y[43];
   assign A[44] = X[44];
   assign B[44] = Y[44];
   assign A[45] = X[45];
   assign B[45] = Y[45];
   assign A[46] = X[46];
   assign B[46] = Y[46];
   assign A[47] = X[47];
   assign B[47] = Y[47];
   assign A[48] = X[48];
   assign B[48] = Y[48];
   assign A[49] = X[49];
   assign B[49] = Y[49];
   assign A[50] = X[50];
   assign B[50] = Y[50];
   assign A[51] = X[51];
   assign B[51] = Y[51];
   assign A[52] = LOGIC0;
   assign B[52] = LOGIC0;
   assign A[53] = LOGIC0;
   assign B[53] = LOGIC0;
   assign A[54] = LOGIC0;
   assign B[54] = LOGIC0;
   assign A[55] = LOGIC0;
   assign B[55] = LOGIC0;
   assign A[56] = LOGIC0;
   assign B[56] = LOGIC0;
   assign A[57] = LOGIC0;
   assign B[57] = LOGIC0;
   assign A[58] = LOGIC0;
   assign B[58] = LOGIC0;
   assign A[59] = LOGIC0;
   assign B[59] = LOGIC0;
   assign A[60] = LOGIC0;
   assign B[60] = LOGIC0;
   assign A[61] = LOGIC0;
   assign B[61] = LOGIC0;
   assign A[62] = LOGIC0;
   assign B[62] = LOGIC0;
   assign A[63] = LOGIC0;
   assign B[63] = LOGIC0;

   assign S[0] = Q[0];
   assign S[1] = Q[1];
   assign S[2] = Q[2];
   assign S[3] = Q[3];
   assign S[4] = Q[4];
   assign S[5] = Q[5];
   assign S[6] = Q[6];
   assign S[7] = Q[7];
   assign S[8] = Q[8];
   assign S[9] = Q[9];
   assign S[10] = Q[10];
   assign S[11] = Q[11];
   assign S[12] = Q[12];
   assign S[13] = Q[13];
   assign S[14] = Q[14];
   assign S[15] = Q[15];
   assign S[16] = Q[16];
   assign S[17] = Q[17];
   assign S[18] = Q[18];
   assign S[19] = Q[19];
   assign S[20] = Q[20];
   assign S[21] = Q[21];
   assign S[22] = Q[22];
   assign S[23] = Q[23];
   assign S[24] = Q[24];
   assign S[25] = Q[25];
   assign S[26] = Q[26];
   assign S[27] = Q[27];
   assign S[28] = Q[28];
   assign S[29] = Q[29];
   assign S[30] = Q[30];
   assign S[31] = Q[31];
   assign S[32] = Q[32];
   assign S[33] = Q[33];
   assign S[34] = Q[34];
   assign S[35] = Q[35];
   assign S[36] = Q[36];
   assign S[37] = Q[37];
   assign S[38] = Q[38];
   assign S[39] = Q[39];
   assign S[40] = Q[40];
   assign S[41] = Q[41];
   assign S[42] = Q[42];
   assign S[43] = Q[43];
   assign S[44] = Q[44];
   assign S[45] = Q[45];
   assign S[46] = Q[46];
   assign S[47] = Q[47];
   assign S[48] = Q[48];
   assign S[49] = Q[49];
   assign S[50] = Q[50];
   assign S[51] = Q[51];
   assign CO_52 = Q[52];
   
endmodule //cla_sub52

///////////////////////////////////////////
// wallypipelinedcore.sv
//
// Written: David_Harris@hmc.edu 9 January 2021
// Modified: 
//
// Purpose: Pipelined RISC-V Processor
// 
// Documentation: RISC-V System on Chip Design (Figure 4.1)
//
// A component of the CORE-V-WALLY configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

import cvw::*;  // global CORE-V-Wally parameters

module wallypipelinedcore #(parameter cvw_t P) (
   input  logic                  clk, reset,
   // Privileged
   input  logic                  MTimerInt, MExtInt, SExtInt, MSwInt,
   input  logic [63:0]           MTIME_CLINT, 
   // Bus Interface
<<<<<<< HEAD
   input  logic [P.AHBW-1:0]       HRDATA,
   input  logic                  HREADY, HRESP,
   output logic                  HCLK, HRESETn,
   output logic [P.PA_BITS-1:0]    HADDR,
   output logic [P.AHBW-1:0]       HWDATA,
   output logic [P.XLEN/8-1:0]     HWSTRB,
=======
   input  logic [`AHBW-1:0]      HRDATA,
   input  logic                  HREADY, HRESP,
   output logic                  HCLK, HRESETn,
   output logic [`PA_BITS-1:0]   HADDR,
   output logic [`AHBW-1:0]      HWDATA,
   output logic [`XLEN/8-1:0]    HWSTRB,
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
   output logic                  HWRITE,
   output logic [2:0]            HSIZE,
   output logic [2:0]            HBURST,
   output logic [3:0]            HPROT,
   output logic [1:0]            HTRANS,
   output logic                  HMASTLOCK
);

  logic                          StallF, StallD, StallE, StallM, StallW;
  logic                          FlushD, FlushE, FlushM, FlushW;
  logic                          RetM;
  logic TrapM;

  //  signals that must connect through DP
  logic                          IntDivE, W64E;
  logic                          CSRReadM, CSRWriteM, PrivilegedM;
  logic [1:0]                    AtomicM;
<<<<<<< HEAD
  logic [P.XLEN-1:0]               ForwardedSrcAE, ForwardedSrcBE;
  logic [P.XLEN-1:0] 			  SrcAM;
  logic [2:0]                    Funct3E;
  logic [31:0]                   InstrD;
  logic [31:0] 					 InstrM, InstrOrigM;
  logic [P.XLEN-1:0]               PCSpillF, PCE, PCLinkE;
  logic [P.XLEN-1:0] 			  PCM;
  logic [P.XLEN-1:0]               CSRReadValW, MDUResultW;
  logic [P.XLEN-1:0]               UnalignedPCNextF, PC2NextF;
  logic [1:0] 					 MemRWM;
  logic 						 InstrValidD, InstrValidE, InstrValidM;
=======
  logic [`XLEN-1:0]              ForwardedSrcAE, ForwardedSrcBE;
  logic [`XLEN-1:0]              SrcAM;
  logic [2:0]                    Funct3E;
  logic [31:0]                   InstrD;
  logic [31:0]                   InstrM, InstrOrigM;
  logic [`XLEN-1:0]              PCSpillF, PCE, PCLinkE;
  logic [`XLEN-1:0]              PCM;
  logic [`XLEN-1:0]              CSRReadValW, MDUResultW;
  logic [`XLEN-1:0]              UnalignedPCNextF, PC2NextF;
  logic [1:0]                    MemRWM;
  logic                          InstrValidD, InstrValidE, InstrValidM;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic                          InstrMisalignedFaultM;
  logic                          IllegalBaseInstrD, IllegalFPUInstrD, IllegalIEUFPUInstrD;
  logic                          InstrPageFaultF, LoadPageFaultM, StoreAmoPageFaultM;
  logic                          LoadMisalignedFaultM, LoadAccessFaultM;
  logic                          StoreAmoMisalignedFaultM, StoreAmoAccessFaultM;
  logic                          InvalidateICacheM, FlushDCacheM;
  logic                          PCSrcE;
  logic                          CSRWriteFenceM;
  logic                          DivBusyE;
  logic                          LoadStallD, StoreStallD, MDUStallD, CSRRdStallD;
  logic                          SquashSCW;

  // floating point unit signals
  logic [2:0]                    FRM_REGW;
  logic [4:0]                    RdE, RdM, RdW;
  logic                          FPUStallD;
  logic                          FWriteIntE;
<<<<<<< HEAD
  logic [P.FLEN-1:0]               FWriteDataM;
  logic [P.XLEN-1:0]               FIntResM;  
  logic [P.XLEN-1:0]              FCvtIntResW; 
=======
  logic [`FLEN-1:0]              FWriteDataM;
  logic [`XLEN-1:0]              FIntResM;  
  logic [`XLEN-1:0]              FCvtIntResW; 
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic                          FCvtIntW; 
  logic                          FDivBusyE;
  logic                          FRegWriteM;
  logic                          FCvtIntStallD;
  logic                          FpLoadStoreM;
  logic [4:0]                    SetFflagsM;
<<<<<<< HEAD
  logic [P.XLEN-1:0]               FIntDivResultW;
=======
  logic [`XLEN-1:0]              FIntDivResultW;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a

  // memory management unit signals
  logic                          ITLBWriteF;
  logic                          ITLBMissF;
<<<<<<< HEAD
  logic [P.XLEN-1:0]               SATP_REGW;
=======
  logic [`XLEN-1:0]              SATP_REGW;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic                          STATUS_MXR, STATUS_SUM, STATUS_MPRV;
  logic [1:0]                    STATUS_MPP, STATUS_FS;
  logic [1:0]                    PrivilegeModeW;
<<<<<<< HEAD
  logic [P.XLEN-1:0]               PTE;
=======
  logic [`XLEN-1:0]              PTE;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic [1:0]                    PageType;
  logic                          sfencevmaM, WFIStallM;
  logic                          SelHPTW;

  // PMA checker signals
<<<<<<< HEAD
  var logic [P.PA_BITS-3:0]           PMPADDR_ARRAY_REGW[P.PMP_ENTRIES-1:0];
  var logic [7:0]                PMPCFG_ARRAY_REGW[P.PMP_ENTRIES-1:0];
=======
  var logic [`PA_BITS-3:0]       PMPADDR_ARRAY_REGW[`PMP_ENTRIES-1:0];
  var logic [7:0]                PMPCFG_ARRAY_REGW[`PMP_ENTRIES-1:0];
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a

  // IMem stalls
  logic                          IFUStallF;
  logic                          LSUStallM;

  // cpu lsu interface
  logic [2:0]                    Funct3M;
<<<<<<< HEAD
  logic [P.XLEN-1:0]               IEUAdrE;
  logic [P.XLEN-1:0]  WriteDataM;
  logic [P.XLEN-1:0]  IEUAdrM;  
  logic [P.LLEN-1:0]               ReadDataW;  
  logic                          CommittedM;

  // AHB ifu interface
  logic [P.PA_BITS-1:0]            IFUHADDR;
=======
  logic [`XLEN-1:0]              IEUAdrE;
  logic [`XLEN-1:0]              WriteDataM;
  logic [`XLEN-1:0]              IEUAdrM;  
  logic [`LLEN-1:0]              ReadDataW;  
  logic                          CommittedM;

  // AHB ifu interface
  logic [`PA_BITS-1:0]           IFUHADDR;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic [2:0]                    IFUHBURST;
  logic [1:0]                    IFUHTRANS;
  logic [2:0]                    IFUHSIZE;
  logic                          IFUHWRITE;
  logic                          IFUHREADY;
  
  // AHB LSU interface
<<<<<<< HEAD
  logic [P.PA_BITS-1:0]            LSUHADDR;
  logic [P.XLEN-1:0]               LSUHWDATA;
  logic [P.XLEN/8-1:0]             LSUHWSTRB;
=======
  logic [`PA_BITS-1:0]           LSUHADDR;
  logic [`XLEN-1:0]              LSUHWDATA;
  logic [`XLEN/8-1:0]            LSUHWSTRB;
>>>>>>> 46e08410112c38dc213a034105f96f6979e1680a
  logic                          LSUHWRITE;
  logic                          LSUHREADY;
  
  logic                          BPWrongE, BPWrongM;
  logic                          BPDirPredWrongM;
  logic                          BTAWrongM;
  logic                          RASPredPCWrongM;
  logic                          IClassWrongM;
  logic [3:0]                    InstrClassM;
  logic                          InstrAccessFaultF, HPTWInstrAccessFaultM;
  logic [2:0]                    LSUHSIZE;
  logic [2:0]                    LSUHBURST;
  logic [1:0]                    LSUHTRANS;
  
  logic                          DCacheMiss;
  logic                          DCacheAccess;
  logic                          ICacheMiss;
  logic                          ICacheAccess;
  logic                          BreakpointFaultM, EcallFaultM;
  logic                          InstrUpdateDAF;
  logic                          BigEndianM;
  logic                          FCvtIntE;
  logic                          CommittedF;
  logic                          BranchD, BranchE, JumpD, JumpE;
  logic                          DCacheStallM, ICacheStallF;
  
  // instruction fetch unit: PC, branch prediction, instruction cache
  ifu ifu(.clk, .reset,
    .StallF, .StallD, .StallE, .StallM, .StallW, .FlushD, .FlushE, .FlushM, .FlushW,
    .InstrValidM, .InstrValidE, .InstrValidD,
    .BranchD, .BranchE, .JumpD, .JumpE, .ICacheStallF,
    // Fetch
    .HRDATA, .PCSpillF, .IFUHADDR, .PC2NextF,
    .IFUStallF, .IFUHBURST, .IFUHTRANS, .IFUHSIZE, .IFUHREADY, .IFUHWRITE,
    .ICacheAccess, .ICacheMiss,
    // Execute
    .PCLinkE, .PCSrcE, .IEUAdrE, .IEUAdrM, .PCE, .BPWrongE,  .BPWrongM, 
    // Mem
    .CommittedF, .UnalignedPCNextF, .InvalidateICacheM, .CSRWriteFenceM,
    .InstrD, .InstrM, .InstrOrigM, .PCM, .InstrClassM, .BPDirPredWrongM,
    .BTAWrongM, .RASPredPCWrongM, .IClassWrongM,
    // Faults out
    .IllegalBaseInstrD, .IllegalFPUInstrD, .InstrPageFaultF, .IllegalIEUFPUInstrD, .InstrMisalignedFaultM,
    // mmu management
    .PrivilegeModeW, .PTE, .PageType, .SATP_REGW, .STATUS_MXR, .STATUS_SUM, .STATUS_MPRV,
    .STATUS_MPP, .ITLBWriteF, .sfencevmaM, .ITLBMissF,
    // pmp/pma (inside mmu) signals. 
    .PMPCFG_ARRAY_REGW,  .PMPADDR_ARRAY_REGW, .InstrAccessFaultF, .InstrUpdateDAF); 
    
  // integer execution unit: integer register file, datapath and controller
  ieu ieu(.clk, .reset,
     // Decode Stage interface
     .InstrD, .IllegalIEUFPUInstrD, .IllegalBaseInstrD,
     // Execute Stage interface
     .PCE, .PCLinkE, .FWriteIntE, .FCvtIntE, .IEUAdrE, .IntDivE, .W64E,
     .Funct3E, .ForwardedSrcAE, .ForwardedSrcBE, 
     // Memory stage interface
     .SquashSCW, // from LSU
     .MemRWM, // read/write control goes to LSU
     .AtomicM, // atomic control goes to LSU
     .WriteDataM, // Write data to LSU
     .Funct3M, // size and signedness to LSU
     .SrcAM, // to privilege and fpu
     .RdE, .RdM, .FIntResM, .FlushDCacheM,
     .BranchD, .BranchE, .JumpD, .JumpE,
     // Writeback stage
     .CSRReadValW, .MDUResultW, .FIntDivResultW, .RdW, .ReadDataW(ReadDataW[P.XLEN-1:0]),
     .InstrValidM, .InstrValidE, .InstrValidD, .FCvtIntResW, .FCvtIntW,
     // hazards
     .StallD, .StallE, .StallM, .StallW, .FlushD, .FlushE, .FlushM, .FlushW,
     .FCvtIntStallD, .LoadStallD, .MDUStallD, .CSRRdStallD, .PCSrcE,
     .CSRReadM, .CSRWriteM, .PrivilegedM, .CSRWriteFenceM, .InvalidateICacheM, .StoreStallD); 

  lsu lsu(
    .clk, .reset, .StallM, .FlushM, .StallW, .FlushW,
    // CPU interface
    .MemRWM, .Funct3M, .Funct7M(InstrM[31:25]), .AtomicM,
    .CommittedM, .DCacheMiss, .DCacheAccess, .SquashSCW,            
    .FpLoadStoreM, .FWriteDataM, .IEUAdrE, .IEUAdrM, .WriteDataM,
    .ReadDataW, .FlushDCacheM,
    // connected to ahb (all stay the same)
    .LSUHADDR,  .HRDATA, .LSUHWDATA, .LSUHWSTRB, .LSUHSIZE, 
    .LSUHBURST, .LSUHTRANS, .LSUHWRITE, .LSUHREADY,
    // connect to csr or privilege and stay the same.
    .PrivilegeModeW, .BigEndianM,          // connects to csr
    .PMPCFG_ARRAY_REGW,     // connects to csr
    .PMPADDR_ARRAY_REGW,    // connects to csr
    // hptw keep i/o
    .SATP_REGW, // from csr
    .STATUS_MXR, // from csr
    .STATUS_SUM,  // from csr
    .STATUS_MPRV,  // from csr            
    .STATUS_MPP,  // from csr      
    .sfencevmaM,                   // connects to privilege
    .DCacheStallM,                  // connects to privilege
    .LoadPageFaultM,   // connects to privilege
    .StoreAmoPageFaultM, // connects to privilege
    .LoadMisalignedFaultM, // connects to privilege
    .LoadAccessFaultM,         // connects to privilege
    .HPTWInstrAccessFaultM,         // connects to privilege
    .StoreAmoMisalignedFaultM, // connects to privilege
    .StoreAmoAccessFaultM,     // connects to privilege
    .InstrUpdateDAF,
    .PCSpillF, .ITLBMissF, .PTE, .PageType, .ITLBWriteF, .SelHPTW,
    .LSUStallM);                    

  if (P.BUS_SUPPORTED) begin : ebu
    ebu ebu(// IFU connections
      .clk, .reset,
      // IFU interface
      .IFUHADDR, .IFUHBURST, .IFUHTRANS, .IFUHREADY, .IFUHSIZE,
      // LSU interface
      .LSUHADDR, .LSUHWDATA, .LSUHWSTRB, .LSUHSIZE, .LSUHBURST,
      .LSUHTRANS, .LSUHWRITE, .LSUHREADY,
      // BUS interface
      .HREADY, .HRESP, .HCLK, .HRESETn,
      .HADDR, .HWDATA, .HWSTRB, .HWRITE, .HSIZE, .HBURST,
      .HPROT, .HTRANS, .HMASTLOCK);
  end

  // global stall and flush control  
  hazard  hzu(
    .BPWrongE, .CSRWriteFenceM, .RetM, .TrapM,
    .LoadStallD, .StoreStallD, .MDUStallD, .CSRRdStallD,
    .LSUStallM, .IFUStallF,
    .FCvtIntStallD, .FPUStallD,
    .DivBusyE, .FDivBusyE,
    .EcallFaultM, .BreakpointFaultM,
    .WFIStallM,
    // Stall & flush outputs
    .StallF, .StallD, .StallE, .StallM, .StallW,
    .FlushD, .FlushE, .FlushM, .FlushW);    

  // privileged unit
  if (P.ZICSR_SUPPORTED) begin:priv
    privileged priv(
      .clk, .reset,
      .FlushD, .FlushE, .FlushM, .FlushW, .StallD, .StallE, .StallM, .StallW,
      .CSRReadM, .CSRWriteM, .SrcAM, .PCM, .PC2NextF,
      .InstrM, .InstrOrigM, .CSRReadValW, .UnalignedPCNextF,
      .RetM, .TrapM, .sfencevmaM, .InvalidateICacheM, .DCacheStallM, .ICacheStallF,
      .InstrValidM, .CommittedM, .CommittedF,
      .FRegWriteM, .LoadStallD, .StoreStallD,
      .BPDirPredWrongM, .BTAWrongM, .BPWrongM,
      .RASPredPCWrongM, .IClassWrongM, .DivBusyE, .FDivBusyE,
      .InstrClassM, .DCacheMiss, .DCacheAccess, .ICacheMiss, .ICacheAccess, .PrivilegedM,
      .InstrPageFaultF, .LoadPageFaultM, .StoreAmoPageFaultM,
      .InstrMisalignedFaultM, .IllegalIEUFPUInstrD, 
      .LoadMisalignedFaultM, .StoreAmoMisalignedFaultM,
      .MTimerInt, .MExtInt, .SExtInt, .MSwInt,
      .MTIME_CLINT, .IEUAdrM, .SetFflagsM,
      .InstrAccessFaultF, .HPTWInstrAccessFaultM, .LoadAccessFaultM, .StoreAmoAccessFaultM, .SelHPTW,
      .PrivilegeModeW, .SATP_REGW,
      .STATUS_MXR, .STATUS_SUM, .STATUS_MPRV, .STATUS_MPP, .STATUS_FS,
      .PMPCFG_ARRAY_REGW, .PMPADDR_ARRAY_REGW, 
      .FRM_REGW,.BreakpointFaultM, .EcallFaultM, .WFIStallM, .BigEndianM);
  end else begin
    assign CSRReadValW = 0;
    assign UnalignedPCNextF = PC2NextF;
    assign RetM = 0;
    assign TrapM = 0;
    assign WFIStallM = 0;
    assign sfencevmaM = 0;
    assign BigEndianM = 0;
  end

  // multiply/divide unit
  if (P.M_SUPPORTED | P.ZMMUL_SUPPORTED) begin:mdu
    mdu mdu(.clk, .reset, .StallM, .StallW, .FlushE, .FlushM, .FlushW,
      .ForwardedSrcAE, .ForwardedSrcBE, 
      .Funct3E, .Funct3M, .IntDivE, .W64E,
      .MDUResultW, .DivBusyE); 
  end else begin // no M instructions supported
    assign MDUResultW = 0; 
    assign DivBusyE = 0;
  end

  // floating point unit
  if (P.F_SUPPORTED) begin:fpu
    fpu fpu(
      .clk, .reset,
      .FRM_REGW, // Rounding mode from CSR
      .InstrD, // instruction from IFU
      .ReadDataW(ReadDataW[P.FLEN-1:0]),// Read data from memory
      .ForwardedSrcAE, // Integer input being processed (from IEU)
      .StallE, .StallM, .StallW, // stall signals from HZU
      .FlushE, .FlushM, .FlushW, // flush signals from HZU
      .RdE, .RdM, .RdW, // which FP register to write to (from IEU)
      .STATUS_FS, // is floating-point enabled?
      .FRegWriteM, // FP register write enable
      .FpLoadStoreM,
      .ForwardedSrcBE, // Integer input for intdiv
      .Funct3E, .Funct3M, .IntDivE, .W64E, // Integer flags and functions
      .FPUStallD, // Stall the decode stage
      .FWriteIntE, .FCvtIntE, // integer register write enable, conversion operation
      .FWriteDataM, // Data to be written to memory
      .FIntResM, // data to be written to integer register
      .FCvtIntResW, // fp -> int conversion result to be stored in int register
      .FCvtIntW,   // fpu result selection
      .FDivBusyE, // Is the divide/sqrt unit busy (stall execute stage)
      .IllegalFPUInstrD, // Is the instruction an illegal fpu instruction
      .SetFflagsM,        // FPU flags (to privileged unit)
      .FIntDivResultW); 
  end else begin // no F_SUPPORTED or D_SUPPORTED; tie outputs low
    assign FPUStallD = 0;
    assign FWriteIntE = 0; 
    assign FCvtIntE = 0;
    assign FIntResM = 0;
    assign FCvtIntW = 0;
    assign FDivBusyE = 0;
    assign IllegalFPUInstrD = 1;
    assign SetFflagsM = 0;
    assign FpLoadStoreM = 0;
  end
  
endmodule

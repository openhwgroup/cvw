///////////////////////////////////////////
// rom1p1r
//
// Written: David_Harris@hmc.edu 8/24/22
//
// Purpose: Single-ported ROM
// 
// A component of the CORE-V-WALLY configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

// This model actually works correctly with vivado.

`include "wally-config.vh"

module rom1p1r #(parameter ADDR_WIDTH = 8,
		 parameter DATA_WIDTH = 32, 
		 parameter PRELOAD_ENABLED = 0)
  (input  logic                  clk,
   input  logic                  ce,
   input  logic [ADDR_WIDTH-1:0] addr,
   output logic [DATA_WIDTH-1:0] dout
);

   // Core Memory
   logic [DATA_WIDTH-1:0] 	 ROM [(2**ADDR_WIDTH)-1:0];
   if (`USE_SRAM == 1 && DATA_WIDTH == 64) begin
      rom1p1r_128x64 rom1 (.CLK(clk), .CEB(~ce), .A(addr[6:0]), .Q(dout));

   end if (`USE_SRAM == 1 && DATA_WIDTH == 32) begin
      rom1p1r_128x32 rom1 (.CLK(clk), .CEB(~ce), .A(addr[6:0]), .Q(dout));      

   end else begin
      always @ (posedge clk) begin
	 if(ce) dout <= ROM[addr];    
      end
   
   // for FPGA, initialize with zero-stage bootloader
   if(PRELOAD_ENABLED) begin
      initial begin
	 /*ROM[0] =  64'h9581819300002197; 
	 ROM[1] =  64'h4281420141014081; 
	 ROM[2] =  64'h4481440143814301; 
	 ROM[3] =  64'h4681460145814501; 
	 ROM[4] =  64'h4881480147814701; 
	 ROM[5] =  64'h4a814a0149814901; 
	 ROM[6] =  64'h4c814c014b814b01; 
	 ROM[7] =  64'h4e814e014d814d01; 
	 ROM[8] =  64'h0110011b4f814f01; 
	 ROM[9] =  64'h059b45011161016e; 
	 ROM[10] = 64'h0004063705fe0010; 
	 ROM[11] = 64'h05a000ef8006061b; 
	 ROM[12] = 64'h0ff003930000100f; 
	 ROM[13] = 64'h4e952e3110060e37; 
	 ROM[14] = 64'hc602829b0053f2b7; 
	 ROM[15] = 64'h2023fe02dfe312fd; 
	 ROM[16] = 64'h829b0053f2b7007e; 
	 ROM[17] = 64'hfe02dfe312fdc602; 
	 ROM[18] = 64'h4de31efd000e2023; 
	 ROM[19] = 64'h059bf1402573fdd0; 
	 ROM[20] = 64'h0000061705e20870; 
	 ROM[21] = 64'h0010029b01260613; 
	 ROM[22] = 64'h11010002806702fe; 
	 ROM[23] = 64'h84b2842ae426e822; 
	 ROM[24] = 64'h892ee04aec064511; 
	 ROM[25] = 64'h06e000ef07e000ef; 
	 ROM[26] = 64'h979334fd02905563; 
	 ROM[27] = 64'h07930177d4930204; 
	 ROM[28] = 64'h4089093394be2004; 
	 ROM[29] = 64'h04138522008905b3; 
	 ROM[30] = 64'h19e3014000ef2004; 
	 ROM[31] = 64'h64a2644260e2fe94; 
	 ROM[32] = 64'h6749808261056902; 
	 ROM[33] = 64'hdfed8b8510472783; 
	 ROM[34] = 64'h2423479110a73823; 
	 ROM[35] = 64'h10472783674910f7; 
	 ROM[36] = 64'h20058693ffed8b89; 
	 ROM[37] = 64'h05a1118737836749; 
	 ROM[38] = 64'hfed59be3fef5bc23; 
	 ROM[39] = 64'h1047278367498082; 
	 ROM[40] = 64'h47858082dfed8b85; 
	 ROM[41] = 64'h40a7853b4015551b;   
	 ROM[42] = 64'h808210a7a02367c9;*/

        ROM[0]  = 64'hc001819300002197;
        ROM[1]  = 64'h4281420141014081;
        ROM[2]  = 64'h4481440143814301;
        ROM[3]  = 64'h4681460145814501;
        ROM[4]  = 64'h4881480147814701;
        ROM[5]  = 64'h4a814a0149814901;
        ROM[6]  = 64'h4c814c014b814b01;
        ROM[7]  = 64'h4e814e014d814d01;
        ROM[8]  = 64'h0110011b4f814f01;
        ROM[9]  = 64'h059b45011161016e;
        ROM[10] = 64'h0004063705fe0010;
        ROM[11] = 64'h1ee000ef8006061b;
        ROM[12] = 64'h0ff003930000100f;
        ROM[13] = 64'h4e952e3110060e37;
        ROM[14] = 64'hc602829b0053f2b7;
        ROM[15] = 64'h2023fe02dfe312fd;
        ROM[16] = 64'h829b0053f2b7007e;
        ROM[17] = 64'hfe02dfe312fdc602;
        ROM[18] = 64'h4de31efd000e2023;
        ROM[19] = 64'h059bf1402573fdd0;
        ROM[20] = 64'h0000061705e20870;
        ROM[21] = 64'h0010029b01260613;
        ROM[22] = 64'h67110002806702fe;
        ROM[23] = 64'h0085179bf0070713;
        ROM[24] = 64'h2781038007138ff9;
        ROM[25] = 64'h7563470508a76a63;
        ROM[26] = 64'h00a71733357902a7;
        ROM[27] = 64'h3285350300001517;
        ROM[28] = 64'h40301537e9598d79;
        ROM[29] = 64'h8d7942250513051a;
        ROM[30] = 64'he35d18177713e149;
        ROM[31] = 64'he79300367713c295;
        ROM[32] = 64'hf330674de3450207;
        ROM[33] = 64'h861bc3701ff00613;
        ROM[34] = 64'h01000637c730fff6;
        ROM[35] = 64'hc35c674dcf10167d;
        ROM[36] = 64'hd31c17fd001007b7;
        ROM[37] = 64'h0007861b5b5cc30c;
        ROM[38] = 64'h674d02072a23dfed;
        ROM[39] = 64'h12634785fffd571c;
        ROM[40] = 64'h80818793471006f6;
        ROM[41] = 64'h4b10474cc3904501;
        ROM[42] = 64'hc7d8c790c3cc4b58;
        ROM[43] = 64'h086007138082e29d;
        ROM[44] = 64'h0a90071300e50c63;
        ROM[45] = 64'h0017e793f8e518e3;
        ROM[46] = 64'hb74901d7e793b761;
        ROM[47] = 64'h674dbfb50197e793;
        ROM[48] = 64'h02072e23dffd5f5c;
        ROM[49] = 64'h8513ff7d569866cd;
        ROM[50] = 64'h053300a03533fff7;
        ROM[51] = 64'h00a7e793808240a0;
        ROM[52] = 64'h71398082557dbfa1;
        ROM[53] = 64'hf8228181ca03e852;
        ROM[54] = 64'hf426fc06ec4ef04a;
        ROM[55] = 64'h008a7a13e05ae456;
        ROM[56] = 64'h1463843289ae892a;
        ROM[57] = 64'h4a8500959993000a;
        ROM[58] = 64'h4549864ac4296b05;
        ROM[59] = 64'h055402630009859b;
        ROM[60] = 64'h008b73630004049b;
        ROM[61] = 64'hecbff0ef86a66485;
        ROM[62] = 64'h45814601468187aa;
        ROM[63] = 64'h0207c8639c054531;
        ROM[64] = 64'h0094979beb7ff0ef;
        ROM[65] = 64'h0205406393811782;
        ROM[66] = 64'h99ba020a1863873e;
        ROM[67] = 64'ha8014501fc4d993e;
        ROM[68] = 64'he93ff0ef45454685;
        ROM[69] = 64'h70e24505fe055ae3;
        ROM[70] = 64'h69e2790274a27442;
        ROM[71] = 64'h61216b026aa26a42;
        ROM[72] = 64'h9301020497138082;
        ROM[73] = 64'hec26f0227179b7f9;
        ROM[74] = 64'he44ef4064705e84a;
        ROM[75] = 64'h842e84aad79867cd;
        ROM[76] = 64'h8b85571c674d8932;
        ROM[77] = 64'hd35c03600793dff5;
        ROM[78] = 64'h571c674d02072423;
        ROM[79] = 64'ha737b00026f3fffd;
        ROM[80] = 64'h27f311f707130007;
        ROM[81] = 64'hfef77de38f95b000;
        ROM[82] = 64'h80018c235b1c674d;
        ROM[83] = 64'he7934f5ccf9d8b89;
        ROM[84] = 64'hb00026f3cf5c0027;
        ROM[85] = 64'h0ff7071305f5e737;
        ROM[86] = 64'h7de38f95b00027f3;
        ROM[87] = 64'h9bf54f5c674dfef7;
        ROM[88] = 64'h9737b00026f3cf5c;
        ROM[89] = 64'h27f367f707130098;
        ROM[90] = 64'hfef77de38f95b000;
        ROM[91] = 64'h4501458146014681;
        ROM[92] = 64'h80818993dd7ff0ef;
        ROM[93] = 64'h0593460146814789;
        ROM[94] = 64'h00f9882345211aa0;
        ROM[95] = 64'ha783e50ddbfff0ef;
        ROM[96] = 64'h17d21aa007130009;
        ROM[97] = 64'h479102e79e6393d1;
        ROM[98] = 64'hf0efa80900f98823;
        ROM[99] = 64'ha78302054663da1f;
        ROM[100]= 64'h46810207cc630009;
        ROM[101]= 64'h0370051345814601;
        ROM[102]= 64'h468187aad87ff0ef;
        ROM[103]= 64'h0513403005b74601;
        ROM[104]= 64'h8522fc07dae30a90;
        ROM[105]= 64'h864a69a270a27402;
        ROM[106]= 64'h614564e2694285a6;
        ROM[107]= 64'hebd18b8583f9b5b9;
        ROM[108]= 64'h4509458146014681;
        ROM[109]= 64'hfc054de3d4fff0ef;
        ROM[110]= 64'h123405b746014681;
        ROM[111]= 64'h44e3d3dff0ef450d;
        ROM[112]= 64'h77c10009a983fc05;
        ROM[113]= 64'h460100f9f9b34681;
        ROM[114]= 64'hd23ff0ef451d85ce;
        ROM[115]= 64'h470567cdfa0547e3;
        ROM[116]= 64'h4737b00026f3d3d8;
        ROM[117]= 64'h27f323f70713000f;
        ROM[118]= 64'hfef77de38f95b000;
        ROM[119]= 64'h46810007ae2367cd;
        ROM[120]= 64'h0370051385ce4601;
        ROM[121]= 64'hf6054de3cefff0ef;
        ROM[122]= 64'h0513458146014681;
        ROM[123]= 64'h44e3cddff0ef0860;
        ROM[124]= 64'h059346014681f605;
        ROM[125]= 64'hccbff0ef45412000;
        ROM[126]= 64'he7930109c783bf99;
        ROM[127]= 64'hb78d00f988230087;
        ROM[128]= 64'h0000000000000000;
        ROM[129]= 64'h0000000000000000;
        ROM[130]= 64'h0000000000000000;
        ROM[131]= 64'h0000000000000000;
        ROM[132]= 64'h0000000000000000;
        ROM[133]= 64'h0000000000000000;
        ROM[134]= 64'h0000000000000000;
        ROM[135]= 64'h0000000000000000;
        ROM[136]= 64'h0000000000000000;
        ROM[137]= 64'h0000000000000000;
        ROM[138]= 64'h0000000000000000;
        ROM[139]= 64'h0000000000000000;
        ROM[140]= 64'h0000000000000000;
        ROM[141]= 64'h0000000000000000;
        ROM[142]= 64'h0000000000000000;
        ROM[143]= 64'h0000000000000000;
        ROM[144]= 64'h0000000000000000;
        ROM[145]= 64'h0000000000000000;
        ROM[146]= 64'h0000000000000000;
        ROM[147]= 64'h0000000000000000;
        ROM[148]= 64'h0000000000000000;
        ROM[149]= 64'h0000000000000000;
        ROM[150]= 64'h0000000000000000;
        ROM[151]= 64'h0000000000000000;
        ROM[152]= 64'h0000000000000000;
        ROM[153]= 64'h0000000000000000;
        ROM[154]= 64'h0000000000000000;
        ROM[155]= 64'h0000000000000000;
        ROM[156]= 64'h0000000000000000;
        ROM[157]= 64'h0000000000000000;
        ROM[158]= 64'h0000000000000000;
        ROM[159]= 64'h0000000000000000;
        ROM[160]= 64'h0000000000000000;
        ROM[161]= 64'h0000000000000000;
        ROM[162]= 64'h0000000000000000;
        ROM[163]= 64'h0000000000000000;
        ROM[164]= 64'h0000000000000000;
        ROM[165]= 64'h0000000000000000;
        ROM[166]= 64'h0000000000000000;
        ROM[167]= 64'h0000000000000000;
        ROM[168]= 64'h0000000000000000;
        ROM[169]= 64'h0000000000000000;
        ROM[170]= 64'h0000000000000000;
        ROM[171]= 64'h0000000000000000;
        ROM[172]= 64'h0000000000000000;
        ROM[173]= 64'h0000000000000000;
        ROM[174]= 64'h0000000000000000;
        ROM[175]= 64'h0000000000000000;
        ROM[176]= 64'h0000000000000000;
        ROM[177]= 64'h0000000000000000;
        ROM[178]= 64'h0000000000000000;
        ROM[179]= 64'h0000000000000000;
        ROM[180]= 64'h0000000000000000;
        ROM[181]= 64'h0000000000000000;
        ROM[182]= 64'h0000000000000000;
        ROM[183]= 64'h0000000000000000;
        ROM[184]= 64'h0000000000000000;
        ROM[185]= 64'h0000000000000000;
        ROM[186]= 64'h0000000000000000;
        ROM[187]= 64'h0000000000000000;
        ROM[188]= 64'h0000000000000000;
        ROM[189]= 64'h0000000000000000;
        ROM[190]= 64'h0000000000000000;
        ROM[191]= 64'h0000000000000000;
        ROM[192]= 64'h0000000000000000;
        ROM[193]= 64'h0000000000000000;
        ROM[194]= 64'h0000000000000000;
        ROM[195]= 64'h0000000000000000;
        ROM[196]= 64'h0000000000000000;
        ROM[197]= 64'h0000000000000000;
        ROM[198]= 64'h0000000000000000;
        ROM[199]= 64'h0000000000000000;
        ROM[200]= 64'h0000000000000000;
        ROM[201]= 64'h0000000000000000;
        ROM[202]= 64'h0000000000000000;
        ROM[203]= 64'h0000000000000000;
        ROM[204]= 64'h0000000000000000;
        ROM[205]= 64'h0000000000000000;
        ROM[206]= 64'h0000000000000000;
        ROM[207]= 64'h0000000000000000;
        ROM[208]= 64'h0000000000000000;
        ROM[209]= 64'h0000000000000000;
        ROM[210]= 64'h0000000000000000;
        ROM[211]= 64'h0000000000000000;
        ROM[212]= 64'h0000000000000000;
        ROM[213]= 64'h0000000000000000;
        ROM[214]= 64'h0000000000000000;
        ROM[215]= 64'h0000000000000000;
        ROM[216]= 64'h0000000000000000;
        ROM[217]= 64'h0000000000000000;
        ROM[218]= 64'h0000000000000000;
        ROM[219]= 64'h0000000000000000;
        ROM[220]= 64'h0000000000000000;
        ROM[221]= 64'h0000000000000000;
        ROM[222]= 64'h0000000000000000;
        ROM[223]= 64'h0000000000000000;
        ROM[224]= 64'h0000000000000000;
        ROM[225]= 64'h0000000000000000;
        ROM[226]= 64'h0000000000000000;
        ROM[227]= 64'h0000000000000000;
        ROM[228]= 64'h0000000000000000;
        ROM[229]= 64'h0000000000000000;
        ROM[230]= 64'h0000000000000000;
        ROM[231]= 64'h0000000000000000;
        ROM[232]= 64'h0000000000000000;
        ROM[233]= 64'h0000000000000000;
        ROM[234]= 64'h0000000000000000;
        ROM[235]= 64'h0000000000000000;
        ROM[236]= 64'h0000000000000000;
        ROM[237]= 64'h0000000000000000;
        ROM[238]= 64'h0000000000000000;
        ROM[239]= 64'h0000000000000000;
        ROM[240]= 64'h0000000000000000;
        ROM[241]= 64'h0000000000000000;
        ROM[242]= 64'h0000000000000000;
        ROM[243]= 64'h0000000000000000;
        ROM[244]= 64'h0000000000000000;
        ROM[245]= 64'h0000000000000000;
        ROM[246]= 64'h0000000000000000;
        ROM[247]= 64'h0000000000000000;
        ROM[248]= 64'h0000000000000000;
        ROM[249]= 64'h0000000000000000;
        ROM[250]= 64'h0000000000000000;
        ROM[251]= 64'h0000000000000000;
        ROM[252]= 64'h0000000000000000;
        ROM[253]= 64'h0000000000000000;
        ROM[254]= 64'h0000000000000000;
        ROM[255]= 64'h0000000000000000;
        ROM[256]= 64'h0000000000000000;
        ROM[257]= 64'h0000000000000000;
        ROM[258]= 64'h0000000000000000;
        ROM[259]= 64'h0000000000000000;
        ROM[260]= 64'h0000000000000000;
        ROM[261]= 64'h0000000000000000;
        ROM[262]= 64'h0000000000000000;
        ROM[263]= 64'h0000000000000000;
        ROM[264]= 64'h0000000000000000;
        ROM[265]= 64'h0000000000000000;
        ROM[266]= 64'h0000000000000000;
        ROM[267]= 64'h0000000000000000;
        ROM[268]= 64'h0000000000000000;
        ROM[269]= 64'h0000000000000000;
        ROM[270]= 64'h0000000000000000;
        ROM[271]= 64'h0000000000000000;
        ROM[272]= 64'h0000000000000000;
        ROM[273]= 64'h0000000000000000;
        ROM[274]= 64'h0000000000000000;
        ROM[275]= 64'h0000000000000000;
        ROM[276]= 64'h0000000000000000;
        ROM[277]= 64'h0000000000000000;
        ROM[278]= 64'h0000000000000000;
        ROM[279]= 64'h0000000000000000;
        ROM[280]= 64'h0000000000000000;
        ROM[281]= 64'h0000000000000000;
        ROM[282]= 64'h0000000000000000;
        ROM[283]= 64'h0000000000000000;
        ROM[284]= 64'h0000000000000000;
        ROM[285]= 64'h0000000000000000;
        ROM[286]= 64'h0000000000000000;
        ROM[287]= 64'h0000000000000000;
        ROM[288]= 64'h0000000000000000;
        ROM[289]= 64'h0000000000000000;
        ROM[290]= 64'h0000000000000000;
        ROM[291]= 64'h0000000000000000;
        ROM[292]= 64'h0000000000000000;
        ROM[293]= 64'h0000000000000000;
        ROM[294]= 64'h0000000000000000;
        ROM[295]= 64'h0000000000000000;
        ROM[296]= 64'h0000000000000000;
        ROM[297]= 64'h0000000000000000;
        ROM[298]= 64'h0000000000000000;
        ROM[299]= 64'h0000000000000000;
        ROM[300]= 64'h0000000000000000;
        ROM[301]= 64'h0000000000000000;
        ROM[302]= 64'h0000000000000000;
        ROM[303]= 64'h0000000000000000;
        ROM[304]= 64'h0000000000000000;
        ROM[305]= 64'h0000000000000000;
        ROM[306]= 64'h0000000000000000;
        ROM[307]= 64'h0000000000000000;
        ROM[308]= 64'h0000000000000000;
        ROM[309]= 64'h0000000000000000;
        ROM[310]= 64'h0000000000000000;
        ROM[311]= 64'h0000000000000000;
        ROM[312]= 64'h0000000000000000;
        ROM[313]= 64'h0000000000000000;
        ROM[314]= 64'h0000000000000000;
        ROM[315]= 64'h0000000000000000;
        ROM[316]= 64'h0000000000000000;
        ROM[317]= 64'h0000000000000000;
        ROM[318]= 64'h0000000000000000;
        ROM[319]= 64'h0000000000000000;
        ROM[320]= 64'h0000000000000000;
        ROM[321]= 64'h0000000000000000;
        ROM[322]= 64'h0000000000000000;
        ROM[323]= 64'h0000000000000000;
        ROM[324]= 64'h0000000000000000;
        ROM[325]= 64'h0000000000000000;
        ROM[326]= 64'h0000000000000000;
        ROM[327]= 64'h0000000000000000;
        ROM[328]= 64'h0000000000000000;
        ROM[329]= 64'h0000000000000000;
        ROM[330]= 64'h0000000000000000;
        ROM[331]= 64'h0000000000000000;
        ROM[332]= 64'h0000000000000000;
        ROM[333]= 64'h0000000000000000;
        ROM[334]= 64'h0000000000000000;
        ROM[335]= 64'h0000000000000000;
        ROM[336]= 64'h0000000000000000;
        ROM[337]= 64'h0000000000000000;
        ROM[338]= 64'h0000000000000000;
        ROM[339]= 64'h0000000000000000;
        ROM[340]= 64'h0000000000000000;
        ROM[341]= 64'h0000000000000000;
        ROM[342]= 64'h0000000000000000;
        ROM[343]= 64'h0000000000000000;
        ROM[344]= 64'h0000000000000000;
        ROM[345]= 64'h0000000000000000;
        ROM[346]= 64'h0000000000000000;
        ROM[347]= 64'h0000000000000000;
        ROM[348]= 64'h0000000000000000;
        ROM[349]= 64'h0000000000000000;
        ROM[350]= 64'h0000000000000000;
        ROM[351]= 64'h0000000000000000;
        ROM[352]= 64'h0000000000000000;
        ROM[353]= 64'h0000000000000000;
        ROM[354]= 64'h0000000000000000;
        ROM[355]= 64'h0000000000000000;
        ROM[356]= 64'h0000000000000000;
        ROM[357]= 64'h0000000000000000;
        ROM[358]= 64'h0000000000000000;
        ROM[359]= 64'h0000000000000000;
        ROM[360]= 64'h0000000000000000;
        ROM[361]= 64'h0000000000000000;
        ROM[362]= 64'h0000000000000000;
        ROM[363]= 64'h0000000000000000;
        ROM[364]= 64'h0000000000000000;
        ROM[365]= 64'h0000000000000000;
        ROM[366]= 64'h0000000000000000;
        ROM[367]= 64'h0000000000000000;
        ROM[368]= 64'h0000000000000000;
        ROM[369]= 64'h0000000000000000;
        ROM[370]= 64'h0000000000000000;
        ROM[371]= 64'h0000000000000000;
        ROM[372]= 64'h0000000000000000;
        ROM[373]= 64'h0000000000000000;
        ROM[374]= 64'h0000000000000000;
        ROM[375]= 64'h0000000000000000;
        ROM[376]= 64'h0000000000000000;
        ROM[377]= 64'h0000000000000000;
        ROM[378]= 64'h0000000000000000;
        ROM[379]= 64'h0000000000000000;
        ROM[380]= 64'h0000000000000000;
        ROM[381]= 64'h0000000000000000;
        ROM[382]= 64'h0000000000000000;
        ROM[383]= 64'h0000000000000000;
        ROM[384]= 64'h0000000000000000;
        ROM[385]= 64'h0000000000000000;
        ROM[386]= 64'h0000000000000000;
        ROM[387]= 64'h0000000000000000;
        ROM[388]= 64'h0000000000000000;
        ROM[389]= 64'h0000000000000000;
        ROM[390]= 64'h0000000000000000;
        ROM[391]= 64'h0000000000000000;
        ROM[392]= 64'h0000000000000000;
        ROM[393]= 64'h0000000000000000;
        ROM[394]= 64'h0000000000000000;
        ROM[395]= 64'h0000000000000000;
        ROM[396]= 64'h0000000000000000;
        ROM[397]= 64'h0000000000000000;
        ROM[398]= 64'h0000000000000000;
        ROM[399]= 64'h0000000000000000;
        ROM[400]= 64'h0000000000000000;
        ROM[401]= 64'h0000000000000000;
        ROM[402]= 64'h0000000000000000;
        ROM[403]= 64'h0000000000000000;
        ROM[404]= 64'h0000000000000000;
        ROM[405]= 64'h0000000000000000;
        ROM[406]= 64'h0000000000000000;
        ROM[407]= 64'h0000000000000000;
        ROM[408]= 64'h0000000000000000;
        ROM[409]= 64'h0000000000000000;
        ROM[410]= 64'h0000000000000000;
        ROM[411]= 64'h0000000000000000;
        ROM[412]= 64'h0000000000000000;
        ROM[413]= 64'h0000000000000000;
        ROM[414]= 64'h0000000000000000;
        ROM[415]= 64'h0000000000000000;
        ROM[416]= 64'h0000000000000000;
        ROM[417]= 64'h0000000000000000;
        ROM[418]= 64'h0000000000000000;
        ROM[419]= 64'h0000000000000000;
        ROM[420]= 64'h0000000000000000;
        ROM[421]= 64'h0000000000000000;
        ROM[422]= 64'h0000000000000000;
        ROM[423]= 64'h0000000000000000;
        ROM[424]= 64'h0000000000000000;
        ROM[425]= 64'h0000000000000000;
        ROM[426]= 64'h0000000000000000;
        ROM[427]= 64'h0000000000000000;
        ROM[428]= 64'h0000000000000000;
        ROM[429]= 64'h0000000000000000;
        ROM[430]= 64'h0000000000000000;
        ROM[431]= 64'h0000000000000000;
        ROM[432]= 64'h0000000000000000;
        ROM[433]= 64'h0000000000000000;
        ROM[434]= 64'h0000000000000000;
        ROM[435]= 64'h0000000000000000;
        ROM[436]= 64'h0000000000000000;
        ROM[437]= 64'h0000000000000000;
        ROM[438]= 64'h0000000000000000;
        ROM[439]= 64'h0000000000000000;
        ROM[440]= 64'h0000000000000000;
        ROM[441]= 64'h0000000000000000;
        ROM[442]= 64'h0000000000000000;
        ROM[443]= 64'h0000000000000000;
        ROM[444]= 64'h0000000000000000;
        ROM[445]= 64'h0000000000000000;
        ROM[446]= 64'h0000000000000000;
        ROM[447]= 64'h0000000000000000;
        ROM[448]= 64'h0000000000000000;
        ROM[449]= 64'h0000000000000000;
        ROM[450]= 64'h0000000000000000;
        ROM[451]= 64'h0000000000000000;
        ROM[452]= 64'h0000000000000000;
        ROM[453]= 64'h0000000000000000;
        ROM[454]= 64'h0000000000000000;
        ROM[455]= 64'h0000000000000000;
        ROM[456]= 64'h0000000000000000;
        ROM[457]= 64'h0000000000000000;
        ROM[458]= 64'h0000000000000000;
        ROM[459]= 64'h0000000000000000;
        ROM[460]= 64'h0000000000000000;
        ROM[461]= 64'h0000000000000000;
        ROM[462]= 64'h0000000000000000;
        ROM[463]= 64'h0000000000000000;
        ROM[464]= 64'h0000000000000000;
        ROM[465]= 64'h0000000000000000;
        ROM[466]= 64'h0000000000000000;
        ROM[467]= 64'h0000000000000000;
        ROM[468]= 64'h0000000000000000;
        ROM[469]= 64'h0000000000000000;
        ROM[470]= 64'h0000000000000000;
        ROM[471]= 64'h0000000000000000;
        ROM[472]= 64'h0000000000000000;
        ROM[473]= 64'h0000000000000000;
        ROM[474]= 64'h0000000000000000;
        ROM[475]= 64'h0000000000000000;
        ROM[476]= 64'h0000000000000000;
        ROM[477]= 64'h0000000000000000;
        ROM[478]= 64'h0000000000000000;
        ROM[479]= 64'h0000000000000000;
        ROM[480]= 64'h0000000000000000;
        ROM[481]= 64'h0000000000000000;
        ROM[482]= 64'h0000000000000000;
        ROM[483]= 64'h0000000000000000;
        ROM[484]= 64'h0000000000000000;
        ROM[485]= 64'h0000000000000000;
        ROM[486]= 64'h0000000000000000;
        ROM[487]= 64'h0000000000000000;
        ROM[488]= 64'h0000000000000000;
        ROM[489]= 64'h0000000000000000;
        ROM[490]= 64'h0000000000000000;
        ROM[491]= 64'h0000000000000000;
        ROM[492]= 64'h0000000000000000;
        ROM[493]= 64'h0000000000000000;
        ROM[494]= 64'h0000000000000000;
        ROM[495]= 64'h0000000000000000;
        ROM[496]= 64'h0000000000000000;
        ROM[497]= 64'h0000000000000000;
        ROM[498]= 64'h0000000000000000;
        ROM[499]= 64'h0000000000000000;
        ROM[500]= 64'h0000000000000000;
        ROM[501]= 64'h0000000000000000;
        ROM[502]= 64'h0000000000000000;
        ROM[503]= 64'h0000000000000000;
        ROM[504]= 64'h0000000000000000;
        ROM[505]= 64'h0000000000000000;
        ROM[506]= 64'h0000000000000000;
        ROM[507]= 64'h0000000000000000;
        ROM[508]= 64'h0000000000000000;
        ROM[509]= 64'h0000000000000000;
        ROM[510]= 64'h0000000000000000;
        ROM[511]= 64'h0000000000000000;
        ROM[512]= 64'h0000000000000000;
        ROM[513]= 64'h0000000000000000;
        ROM[514]= 64'h0000000000000000;
        ROM[515]= 64'h0000000000000000;
        ROM[516]= 64'h0000000000000000;
        ROM[517]= 64'h0000000000000000;
        ROM[518]= 64'h0000000000000000;
        ROM[519]= 64'h0000000000000000;
        ROM[520]= 64'h0000000000000000;
        ROM[521]= 64'h0000000000000000;
        ROM[522]= 64'h0000000000000000;
        ROM[523]= 64'h0000000000000000;
        ROM[524]= 64'h0000000000000000;
        ROM[525]= 64'h0000000000000000;
        ROM[526]= 64'h0000000000000000;
        ROM[527]= 64'h0000000000000000;
        ROM[528]= 64'h0000000000000000;
        ROM[529]= 64'h0000000000000000;
        ROM[530]= 64'h0000000000000000;
        ROM[531]= 64'h0000000000000000;
        ROM[532]= 64'h0000000000000000;
        ROM[533]= 64'h0000000000000000;
        ROM[534]= 64'h0000000000000000;
        ROM[535]= 64'h0000000000000000;
        ROM[536]= 64'h0000000000000000;
        ROM[537]= 64'h0000000000000000;
        ROM[538]= 64'h0000000000000000;
        ROM[539]= 64'h0000000000000000;
        ROM[540]= 64'h0000000000000000;
        ROM[541]= 64'h0000000000000000;
        ROM[542]= 64'h0000000000000000;
        ROM[543]= 64'h0000000000000000;
        ROM[544]= 64'h0000000000000000;
        ROM[545]= 64'h0000000000000000;
        ROM[546]= 64'h0000000000000000;
        ROM[547]= 64'h0000000000000000;
        ROM[548]= 64'h0000000000000000;
        ROM[549]= 64'h0000000000000000;
        ROM[550]= 64'h0000000000000000;
        ROM[551]= 64'h0000000000000000;
        ROM[552]= 64'h0000000000000000;
        ROM[553]= 64'h0000000000000000;
        ROM[554]= 64'h0000000000000000;
        ROM[555]= 64'h0000000000000000;
        ROM[556]= 64'h0000000000000000;
        ROM[557]= 64'h0000000000000000;
        ROM[558]= 64'h0000000000000000;
        ROM[559]= 64'h0000000000000000;
        ROM[560]= 64'h0000000000000000;
        ROM[561]= 64'h0000000000000000;
        ROM[562]= 64'h0000000000000000;
        ROM[563]= 64'h0000000000000000;
        ROM[564]= 64'h0000000000000000;
        ROM[565]= 64'h0000000000000000;
        ROM[566]= 64'h0000000000000000;
        ROM[567]= 64'h0000000000000000;
        ROM[568]= 64'h0000000000000000;
        ROM[569]= 64'h0000000000000000;
        ROM[570]= 64'h0000000000000000;
        ROM[571]= 64'h0000000000000000;
        ROM[572]= 64'h0000000000000000;
        ROM[573]= 64'h0000000000000000;
        ROM[574]= 64'h0000000000000000;
        ROM[575]= 64'h0000000000000000;
        ROM[576]= 64'h0000000000000000;
        ROM[577]= 64'h0000000000000000;
        ROM[578]= 64'h0000000000000000;
        ROM[579]= 64'h0000000000000000;
        ROM[580]= 64'h0000000000000000;
        ROM[581]= 64'h0000000000000000;
        ROM[582]= 64'h0000000000000000;
        ROM[583]= 64'h0000000000000000;
        ROM[584]= 64'h0000000000000000;
        ROM[585]= 64'h0000000000000000;
        ROM[586]= 64'h0000000000000000;
        ROM[587]= 64'h0000000000000000;
        ROM[588]= 64'h0000000000000000;
        ROM[589]= 64'h0000000000000000;
        ROM[590]= 64'h0000000000000000;
        ROM[591]= 64'h0000000000000000;
        ROM[592]= 64'h0000000000000000;
        ROM[593]= 64'h0000000000000000;
        ROM[594]= 64'h0000000000000000;
        ROM[595]= 64'h0000000000000000;
        ROM[596]= 64'h0000000000000000;
        ROM[597]= 64'h0000000000000000;
        ROM[598]= 64'h0000000000000000;
        ROM[599]= 64'h0000000000000000;
        ROM[600]= 64'h0000000000000000;
        ROM[601]= 64'h0000000000000000;
        ROM[602]= 64'h0000000000000000;
        ROM[603]= 64'h0000000000000000;
        ROM[604]= 64'h0000000000000000;
        ROM[605]= 64'h0000000000000000;
        ROM[606]= 64'h0000000000000000;
        ROM[607]= 64'h0000000000000000;
        ROM[608]= 64'h0000000000000000;
        ROM[609]= 64'h0000000000000000;
        ROM[610]= 64'h0000000000000000;
        ROM[611]= 64'h0000000000000000;
        ROM[612]= 64'h0000000000000000;
        ROM[613]= 64'h0000000000000000;
        ROM[614]= 64'h0000000000000000;
        ROM[615]= 64'h0000000000000000;
        ROM[616]= 64'h0000000000000000;
        ROM[617]= 64'h0000000000000000;
        ROM[618]= 64'h0000000000000000;
        ROM[619]= 64'h0000000000000000;
        ROM[620]= 64'h0000000000000000;
        ROM[621]= 64'h0000000000000000;
        ROM[622]= 64'h0000000000000000;
        ROM[623]= 64'h0000000000000000;
        ROM[624]= 64'h0000000000000000;
        ROM[625]= 64'h0000000000000000;
        ROM[626]= 64'h0000000000000000;
        ROM[627]= 64'h0000000000000000;
        ROM[628]= 64'h0000000000000000;
        ROM[629]= 64'h0000000000000000;
        ROM[630]= 64'h0000000000000000;
        ROM[631]= 64'h0000000000000000;
        ROM[632]= 64'h0000000000000000;
        ROM[633]= 64'h0000000000000000;
        ROM[634]= 64'h0000000000000000;
        ROM[635]= 64'h0000000000000000;
        ROM[636]= 64'h0000000000000000;
        ROM[637]= 64'h0000000000000000;
        ROM[638]= 64'h0000000000000000;
        ROM[639]= 64'h0000000000000000;
        ROM[640]= 64'h00600100d2e3ca40;
      end 
    end 
  end 

endmodule 

///////////////////////////////////////////
// postprocess.sv
//
// Written: kekim@hmc.edu
// Modified: 19 May 2023
//
// Purpose: Post-Processing: normalization, rounding, sign, flags, special cases
// 
// Documentation: RISC-V System on Chip Design Chapter 13
//
// A component of the CORE-V-WALLY configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`include "wally-config.vh"

module divremsqrtpostprocess (
  // general signals
  input logic                             Xs, Ys,     // input signs
  input logic  [`NF:0]                    Xm, Ym,     // input mantissas
  input logic  [2:0]                      Frm,        // rounding mode 000 = rount to nearest, ties to even   001 = round twords zero  010 = round down  011 = round up  100 = round to nearest, ties to max magnitude
  input logic  [`FMTBITS-1:0]             Fmt,        // precision 1 = double 0 = single
  input logic  [2:0]                      OpCtrl,     // choose which opperation (look below for values)
  input logic                             XZero, YZero,        // inputs are zero
  input logic                             XInf, YInf,          // inputs are infinity
  input logic                             XNaN, YNaN,          // inputs are NaN
  input logic                             XSNaN, YSNaN,        // inputs are signaling NaNs
  input logic  [1:0]                      PostProcSel,         // select result to be written to fp register
  //fma signals
  //divide signals
  input logic                             DivSticky,  // divider sticky bit
  input logic  [`NE+1:0]                  DivQe,      // divsqrt exponent
  input logic  [`DIVb:0]                  DivQm,      // divsqrt significand
  // final results
  output logic [`FLEN-1:0]                PostProcRes,// postprocessor final result
  output logic [4:0]                      PostProcFlg // postprocesser flags
  );
  
  // general signals
  logic                       Rs;         // result sign
  logic [`NF-1:0]             Rf;         // Result fraction
  logic [`NE-1:0]             Re;         // Result exponent
  logic                       Ms;         // norMalized sign
  logic [`CORRSHIFTSZ-1:0]    Mf;         // norMalized fraction
  logic [`NE+1:0]             Me;         // normalized exponent
  logic [`NE+1:0]             FullRe;     // Re with bits to determine sign and overflow
  logic                       UfPlus1;    // do you add one (for determining underflow flag)
  logic [`LOGNORMSHIFTSZ-1:0] ShiftAmt;   // normalization shift amount
  logic [`NORMSHIFTSZ-1:0]    ShiftIn;    // input to normalization shift
  logic [`NORMSHIFTSZ-1:0]    Shifted;    // the ouput of the normalized shifter (before shift correction)
  logic                       Plus1;      // add one to the final result?
  logic                       Overflow;   // overflow flag used to select results
  logic                       Invalid;    // invalid flag used to select results
  logic                       Guard, Round, Sticky; // bits needed to determine rounding
  logic [`FMTBITS-1:0]        OutFmt;     // output format
  // division singals
  logic [`LOGNORMSHIFTSZ-1:0] DivShiftAmt;        // divsqrt shif amount
  logic [`NORMSHIFTSZ-1:0]    DivShiftIn;         // divsqrt shift input
  logic [`NE+1:0]             Qe;                 // divsqrt corrected exponent after corretion shift
  logic                       DivByZero;          // divide by zero flag
  logic                       DivResSubnorm;      // is the divsqrt result subnormal
  logic                       DivSubnormShiftPos; // is the divsqrt subnorm shift amout positive (not underflowed)
  // conversion signals
  logic [`CVTLEN+`NF:0]       CvtShiftIn;         // number to be shifted for converter
  logic [1:0]                 CvtNegResMsbs;      // most significant bits of possibly negated int result
  logic [`XLEN+1:0]           CvtNegRes;          // possibly negated integer result
  logic                       CvtResUf;           // did the convert result underflow
  logic                       IntInvalid;         // invalid integer flag
  // readability signals
  logic                       Mult;       // multiply opperation
  logic                       Sqrt;       // is the divsqrt opperation sqrt
  logic                       Int64;      // is the integer 64 bits?
  logic                       Signed;     // is the opperation with a signed integer?
  logic                       IntToFp;    // is the opperation an int->fp conversion?
  logic                       CvtOp;      // convertion opperation
  logic                       DivOp;      // divider opperation
  logic                       InfIn;      // are any of the inputs infinity
  logic                       NaNIn;      // are any of the inputs NaN

  // signals to help readability
  //assign Signed =  OpCtrl[0];
  //assign Int64 =   OpCtrl[1];
  //assign IntToFp = OpCtrl[2];
  //assign Mult = OpCtrl[2]&~OpCtrl[1]&~OpCtrl[0];
  //assign CvtOp = (PostProcSel == 2'b00);
  //assign FmaOp = (PostProcSel == 2'b10);
  assign DivOp = (PostProcSel == 2'b01);
  assign Sqrt =  OpCtrl[0];

  // is there an input of infinity or NaN being used
  assign InfIn = XInf|YInf;
  assign NaNIn = XNaN|YNaN;

  // choose the ouptut format depending on the opperation
  //      - fp -> fp: OpCtrl contains the percision of the output
  //      - otherwise: Fmt contains the percision of the output
  if (`FPSIZES == 2) 
      //assign OutFmt = IntToFp|~CvtOp ? Fmt : (OpCtrl[1:0] == `FMT); 
      assign OutFmt = Fmt;
  else if (`FPSIZES == 3 | `FPSIZES == 4) 
      //assign OutFmt = IntToFp|~CvtOp ? Fmt : OpCtrl[1:0]; 
      assign OutFmt = Fmt;

  ///////////////////////////////////////////////////////////////////////////////
  // Normalization
  ///////////////////////////////////////////////////////////////////////////////

  // final claulations before shifting
  /*cvtshiftcalc cvtshiftcalc(.ToInt, .CvtCe, .CvtResSubnormUf, .Xm, .CvtLzcIn,  
      .XZero, .IntToFp, .OutFmt, .CvtResUf, .CvtShiftIn);*/

  divshiftcalc divshiftcalc(.DivQe, .DivQm, .DivResSubnorm, .DivSubnormShiftPos, .DivShiftAmt, .DivShiftIn);

  assign ShiftAmt = DivShiftAmt;
  assign ShiftIn = DivShiftIn;
  
  // main normalization shift
  normshift normshift (.ShiftIn, .ShiftAmt, .Shifted);

  // correct for LZA/divsqrt error
  divremsqrtshiftcorrection shiftcorrection(.DivResSubnorm, .DivSubnormShiftPos, .DivOp, .DivQe, .Qe, .Shifted, .Mf);

  ///////////////////////////////////////////////////////////////////////////////
  // Rounding
  ///////////////////////////////////////////////////////////////////////////////

  // round to nearest even
  // round to zero
  // round to -infinity
  // round to infinity
  // round to nearest max magnitude

  // calulate result sign used in rounding unit
  divremsqrtroundsign roundsign( .DivOp, .Sqrt, .Xs, .Ys, Ms);

  divremsqrtround round(.OutFmt, .Frm, .Plus1, .Qe,
      .Ms, .Mf, .DivSticky, .DivOp, .UfPlus1, .FullRe, .Rf, .Re, .Sticky, .Round, .Guard, .Me);

  ///////////////////////////////////////////////////////////////////////////////
  // Sign calculation
  ///////////////////////////////////////////////////////////////////////////////

  /*resultsign resultsign(.Frm, .FmaPs, .FmaAs, .Round, .Sticky, .Guard,
      .FmaOp, .ZInf, .InfIn, .FmaSZero, .Mult, .Ms, .Rs);*/
  assign Rs = Ms;

  ///////////////////////////////////////////////////////////////////////////////
  // Flags
  ///////////////////////////////////////////////////////////////////////////////

  divremsqrtflags flags(.XSNaN, .YSNaN, .XInf, .YInf, .InfIn, .XZero, .YZero, 
              .Xs, .OutFmt, .Sqrt,
              .NaNIn, .Round, .DivByZero,
              .Guard, .Sticky, .UfPlus1,.DivOp, .FullRe, .Plus1,
              .Me, .Invalid, .Overflow, .PostProcFlg);

  ///////////////////////////////////////////////////////////////////////////////
  // Select the result
  ///////////////////////////////////////////////////////////////////////////////

  //negateintres negateintres(.Xs, .Shifted, .Signed, .Int64, .Plus1, .CvtNegResMsbs, .CvtNegRes);

  divremsqrtspecialcase specialcase(.Xs, .Xm, .Ym, .XZero, 
      .Frm, .OutFmt, .XNaN, .YNaN,  
      .NaNIn, .Plus1, .Invalid, .Overflow, .InfIn,
      .XInf, .YInf, .DivOp, .DivByZero, .FullRe, .Rs, .Re, .Rf, .PostProcRes );

endmodule

`include "wally-config.vh"
`define DIVLEN ((`NF<(`XLEN)) ? (`XLEN) : `NF)

module qsel4 (
	input logic [`DIVLEN+3:0] D,
	input logic [`DIVLEN+3:0] WS, WC,
	output logic [3:0] q
);
	logic [6:0] Wmsbs;
	logic [7:0] PreWmsbs;
	logic [2:0] Dmsbs;
	assign PreWmsbs = WC[`DIVLEN+3:`DIVLEN-4] + WS[`DIVLEN+3:`DIVLEN-4];
	assign Wmsbs = PreWmsbs[7:1];
        assign Dmsbs = D[`DIVLEN-1:`DIVLEN-3];
	// D = 0001.xxx...
	// Dmsbs = |   |
    // W =      xxxx.xxx...
	// Wmsbs = |        |

	always_comb
	case({Dmsbs,Wmsbs})
		10'b000_0000000: q = 4'b0000;
		10'b000_0000001: q = 4'b0000;
		10'b000_0000010: q = 4'b0000;
		10'b000_0000011: q = 4'b0000;
		10'b000_0000100: q = 4'b0100;
		10'b000_0000101: q = 4'b0100;
		10'b000_0000110: q = 4'b0100;
		10'b000_0000111: q = 4'b0100;
		10'b000_0001000: q = 4'b0100;
		10'b000_0001001: q = 4'b0100;
		10'b000_0001010: q = 4'b0100;
		10'b000_0001011: q = 4'b0100;
		10'b000_0001100: q = 4'b1000;
		10'b000_0001101: q = 4'b1000;
		10'b000_0001110: q = 4'b1000;
		10'b000_0001111: q = 4'b1000;
		10'b000_0010000: q = 4'b1000;
		10'b000_0010001: q = 4'b1000;
		10'b000_0010010: q = 4'b1000;
		10'b000_0010011: q = 4'b1000;
		10'b000_0010100: q = 4'b1000;
		10'b000_0010101: q = 4'b1000;
		10'b000_0010110: q = 4'b1000;
		10'b000_0010111: q = 4'b1000;
		10'b000_0011000: q = 4'b1000;
		10'b000_0011001: q = 4'b1000;
		10'b000_0011010: q = 4'b1000;
		10'b000_0011011: q = 4'b1000;
		10'b000_0011100: q = 4'b1000;
		10'b000_0011101: q = 4'b1000;
		10'b000_0011110: q = 4'b1000;
		10'b000_0011111: q = 4'b1000;
		10'b000_0100000: q = 4'b1000;
		10'b000_0100001: q = 4'b1000;
		10'b000_0100010: q = 4'b1000;
		10'b000_0100011: q = 4'b1000;
		10'b000_0100100: q = 4'b1000;
		10'b000_0100101: q = 4'b1000;
		10'b000_0100110: q = 4'b1000;
		10'b000_0100111: q = 4'b1000;
		10'b000_0101000: q = 4'b1000;
		10'b000_0101001: q = 4'b1000;
		10'b000_0101010: q = 4'b1000;
		10'b000_0101011: q = 4'b1000;
		10'b000_0101100: q = 4'b1000;
		10'b000_0101101: q = 4'b1000;
		10'b000_0101110: q = 4'b1000;
		10'b000_0101111: q = 4'b1000;
		10'b000_0110000: q = 4'b1000;
		10'b000_0110001: q = 4'b1000;
		10'b000_0110010: q = 4'b1000;
		10'b000_0110011: q = 4'b1000;
		10'b000_0110100: q = 4'b1000;
		10'b000_0110101: q = 4'b1000;
		10'b000_0110110: q = 4'b1000;
		10'b000_0110111: q = 4'b1000;
		10'b000_0111000: q = 4'b1000;
		10'b000_0111001: q = 4'b1000;
		10'b000_0111010: q = 4'b1000;
		10'b000_0111011: q = 4'b1000;
		10'b000_0111100: q = 4'b1000;
		10'b000_0111101: q = 4'b1000;
		10'b000_0111110: q = 4'b1000;
		10'b000_0111111: q = 4'b1000;
		10'b000_1000000: q = 4'b0001;
		10'b000_1000001: q = 4'b0001;
		10'b000_1000010: q = 4'b0001;
		10'b000_1000011: q = 4'b0001;
		10'b000_1000100: q = 4'b0001;
		10'b000_1000101: q = 4'b0001;
		10'b000_1000110: q = 4'b0001;
		10'b000_1000111: q = 4'b0001;
		10'b000_1001000: q = 4'b0001;
		10'b000_1001001: q = 4'b0001;
		10'b000_1001010: q = 4'b0001;
		10'b000_1001011: q = 4'b0001;
		10'b000_1001100: q = 4'b0001;
		10'b000_1001101: q = 4'b0001;
		10'b000_1001110: q = 4'b0001;
		10'b000_1001111: q = 4'b0001;
		10'b000_1010000: q = 4'b0001;
		10'b000_1010001: q = 4'b0001;
		10'b000_1010010: q = 4'b0001;
		10'b000_1010011: q = 4'b0001;
		10'b000_1010100: q = 4'b0001;
		10'b000_1010101: q = 4'b0001;
		10'b000_1010110: q = 4'b0001;
		10'b000_1010111: q = 4'b0001;
		10'b000_1011000: q = 4'b0001;
		10'b000_1011001: q = 4'b0001;
		10'b000_1011010: q = 4'b0001;
		10'b000_1011011: q = 4'b0001;
		10'b000_1011100: q = 4'b0001;
		10'b000_1011101: q = 4'b0001;
		10'b000_1011110: q = 4'b0001;
		10'b000_1011111: q = 4'b0001;
		10'b000_1100000: q = 4'b0001;
		10'b000_1100001: q = 4'b0001;
		10'b000_1100010: q = 4'b0001;
		10'b000_1100011: q = 4'b0001;
		10'b000_1100100: q = 4'b0001;
		10'b000_1100101: q = 4'b0001;
		10'b000_1100110: q = 4'b0001;
		10'b000_1100111: q = 4'b0001;
		10'b000_1101000: q = 4'b0001;
		10'b000_1101001: q = 4'b0001;
		10'b000_1101010: q = 4'b0001;
		10'b000_1101011: q = 4'b0001;
		10'b000_1101100: q = 4'b0001;
		10'b000_1101101: q = 4'b0001;
		10'b000_1101110: q = 4'b0001;
		10'b000_1101111: q = 4'b0001;
		10'b000_1110000: q = 4'b0001;
		10'b000_1110001: q = 4'b0001;
		10'b000_1110010: q = 4'b0001;
		10'b000_1110011: q = 4'b0010;
		10'b000_1110100: q = 4'b0010;
		10'b000_1110101: q = 4'b0010;
		10'b000_1110110: q = 4'b0010;
		10'b000_1110111: q = 4'b0010;
		10'b000_1111000: q = 4'b0010;
		10'b000_1111001: q = 4'b0010;
		10'b000_1111010: q = 4'b0010;
		10'b000_1111011: q = 4'b0010;
		10'b000_1111100: q = 4'b0000;
		10'b000_1111101: q = 4'b0000;
		10'b000_1111110: q = 4'b0000;
		10'b000_1111111: q = 4'b0000;
		10'b001_0000000: q = 4'b0000;
		10'b001_0000001: q = 4'b0000;
		10'b001_0000010: q = 4'b0000;
		10'b001_0000011: q = 4'b0000;
		10'b001_0000100: q = 4'b0100;
		10'b001_0000101: q = 4'b0100;
		10'b001_0000110: q = 4'b0100;
		10'b001_0000111: q = 4'b0100;
		10'b001_0001000: q = 4'b0100;
		10'b001_0001001: q = 4'b0100;
		10'b001_0001010: q = 4'b0100;
		10'b001_0001011: q = 4'b0100;
		10'b001_0001100: q = 4'b0100;
		10'b001_0001101: q = 4'b0100;
		10'b001_0001110: q = 4'b1000;
		10'b001_0001111: q = 4'b1000;
		10'b001_0010000: q = 4'b1000;
		10'b001_0010001: q = 4'b1000;
		10'b001_0010010: q = 4'b1000;
		10'b001_0010011: q = 4'b1000;
		10'b001_0010100: q = 4'b1000;
		10'b001_0010101: q = 4'b1000;
		10'b001_0010110: q = 4'b1000;
		10'b001_0010111: q = 4'b1000;
		10'b001_0011000: q = 4'b1000;
		10'b001_0011001: q = 4'b1000;
		10'b001_0011010: q = 4'b1000;
		10'b001_0011011: q = 4'b1000;
		10'b001_0011100: q = 4'b1000;
		10'b001_0011101: q = 4'b1000;
		10'b001_0011110: q = 4'b1000;
		10'b001_0011111: q = 4'b1000;
		10'b001_0100000: q = 4'b1000;
		10'b001_0100001: q = 4'b1000;
		10'b001_0100010: q = 4'b1000;
		10'b001_0100011: q = 4'b1000;
		10'b001_0100100: q = 4'b1000;
		10'b001_0100101: q = 4'b1000;
		10'b001_0100110: q = 4'b1000;
		10'b001_0100111: q = 4'b1000;
		10'b001_0101000: q = 4'b1000;
		10'b001_0101001: q = 4'b1000;
		10'b001_0101010: q = 4'b1000;
		10'b001_0101011: q = 4'b1000;
		10'b001_0101100: q = 4'b1000;
		10'b001_0101101: q = 4'b1000;
		10'b001_0101110: q = 4'b1000;
		10'b001_0101111: q = 4'b1000;
		10'b001_0110000: q = 4'b1000;
		10'b001_0110001: q = 4'b1000;
		10'b001_0110010: q = 4'b1000;
		10'b001_0110011: q = 4'b1000;
		10'b001_0110100: q = 4'b1000;
		10'b001_0110101: q = 4'b1000;
		10'b001_0110110: q = 4'b1000;
		10'b001_0110111: q = 4'b1000;
		10'b001_0111000: q = 4'b1000;
		10'b001_0111001: q = 4'b1000;
		10'b001_0111010: q = 4'b1000;
		10'b001_0111011: q = 4'b1000;
		10'b001_0111100: q = 4'b1000;
		10'b001_0111101: q = 4'b1000;
		10'b001_0111110: q = 4'b1000;
		10'b001_0111111: q = 4'b1000;
		10'b001_1000000: q = 4'b0001;
		10'b001_1000001: q = 4'b0001;
		10'b001_1000010: q = 4'b0001;
		10'b001_1000011: q = 4'b0001;
		10'b001_1000100: q = 4'b0001;
		10'b001_1000101: q = 4'b0001;
		10'b001_1000110: q = 4'b0001;
		10'b001_1000111: q = 4'b0001;
		10'b001_1001000: q = 4'b0001;
		10'b001_1001001: q = 4'b0001;
		10'b001_1001010: q = 4'b0001;
		10'b001_1001011: q = 4'b0001;
		10'b001_1001100: q = 4'b0001;
		10'b001_1001101: q = 4'b0001;
		10'b001_1001110: q = 4'b0001;
		10'b001_1001111: q = 4'b0001;
		10'b001_1010000: q = 4'b0001;
		10'b001_1010001: q = 4'b0001;
		10'b001_1010010: q = 4'b0001;
		10'b001_1010011: q = 4'b0001;
		10'b001_1010100: q = 4'b0001;
		10'b001_1010101: q = 4'b0001;
		10'b001_1010110: q = 4'b0001;
		10'b001_1010111: q = 4'b0001;
		10'b001_1011000: q = 4'b0001;
		10'b001_1011001: q = 4'b0001;
		10'b001_1011010: q = 4'b0001;
		10'b001_1011011: q = 4'b0001;
		10'b001_1011100: q = 4'b0001;
		10'b001_1011101: q = 4'b0001;
		10'b001_1011110: q = 4'b0001;
		10'b001_1011111: q = 4'b0001;
		10'b001_1100000: q = 4'b0001;
		10'b001_1100001: q = 4'b0001;
		10'b001_1100010: q = 4'b0001;
		10'b001_1100011: q = 4'b0001;
		10'b001_1100100: q = 4'b0001;
		10'b001_1100101: q = 4'b0001;
		10'b001_1100110: q = 4'b0001;
		10'b001_1100111: q = 4'b0001;
		10'b001_1101000: q = 4'b0001;
		10'b001_1101001: q = 4'b0001;
		10'b001_1101010: q = 4'b0001;
		10'b001_1101011: q = 4'b0001;
		10'b001_1101100: q = 4'b0001;
		10'b001_1101101: q = 4'b0001;
		10'b001_1101110: q = 4'b0001;
		10'b001_1101111: q = 4'b0001;
		10'b001_1110000: q = 4'b0001;
		10'b001_1110001: q = 4'b0010;
		10'b001_1110010: q = 4'b0010;
		10'b001_1110011: q = 4'b0010;
		10'b001_1110100: q = 4'b0010;
		10'b001_1110101: q = 4'b0010;
		10'b001_1110110: q = 4'b0010;
		10'b001_1110111: q = 4'b0010;
		10'b001_1111000: q = 4'b0010;
		10'b001_1111001: q = 4'b0010;
		10'b001_1111010: q = 4'b0000;
		10'b001_1111011: q = 4'b0000;
		10'b001_1111100: q = 4'b0000;
		10'b001_1111101: q = 4'b0000;
		10'b001_1111110: q = 4'b0000;
		10'b001_1111111: q = 4'b0000;
		10'b010_0000000: q = 4'b0000;
		10'b010_0000001: q = 4'b0000;
		10'b010_0000010: q = 4'b0000;
		10'b010_0000011: q = 4'b0000;
		10'b010_0000100: q = 4'b0100;
		10'b010_0000101: q = 4'b0100;
		10'b010_0000110: q = 4'b0100;
		10'b010_0000111: q = 4'b0100;
		10'b010_0001000: q = 4'b0100;
		10'b010_0001001: q = 4'b0100;
		10'b010_0001010: q = 4'b0100;
		10'b010_0001011: q = 4'b0100;
		10'b010_0001100: q = 4'b0100;
		10'b010_0001101: q = 4'b0100;
		10'b010_0001110: q = 4'b0100;
		10'b010_0001111: q = 4'b1000;
		10'b010_0010000: q = 4'b1000;
		10'b010_0010001: q = 4'b1000;
		10'b010_0010010: q = 4'b1000;
		10'b010_0010011: q = 4'b1000;
		10'b010_0010100: q = 4'b1000;
		10'b010_0010101: q = 4'b1000;
		10'b010_0010110: q = 4'b1000;
		10'b010_0010111: q = 4'b1000;
		10'b010_0011000: q = 4'b1000;
		10'b010_0011001: q = 4'b1000;
		10'b010_0011010: q = 4'b1000;
		10'b010_0011011: q = 4'b1000;
		10'b010_0011100: q = 4'b1000;
		10'b010_0011101: q = 4'b1000;
		10'b010_0011110: q = 4'b1000;
		10'b010_0011111: q = 4'b1000;
		10'b010_0100000: q = 4'b1000;
		10'b010_0100001: q = 4'b1000;
		10'b010_0100010: q = 4'b1000;
		10'b010_0100011: q = 4'b1000;
		10'b010_0100100: q = 4'b1000;
		10'b010_0100101: q = 4'b1000;
		10'b010_0100110: q = 4'b1000;
		10'b010_0100111: q = 4'b1000;
		10'b010_0101000: q = 4'b1000;
		10'b010_0101001: q = 4'b1000;
		10'b010_0101010: q = 4'b1000;
		10'b010_0101011: q = 4'b1000;
		10'b010_0101100: q = 4'b1000;
		10'b010_0101101: q = 4'b1000;
		10'b010_0101110: q = 4'b1000;
		10'b010_0101111: q = 4'b1000;
		10'b010_0110000: q = 4'b1000;
		10'b010_0110001: q = 4'b1000;
		10'b010_0110010: q = 4'b1000;
		10'b010_0110011: q = 4'b1000;
		10'b010_0110100: q = 4'b1000;
		10'b010_0110101: q = 4'b1000;
		10'b010_0110110: q = 4'b1000;
		10'b010_0110111: q = 4'b1000;
		10'b010_0111000: q = 4'b1000;
		10'b010_0111001: q = 4'b1000;
		10'b010_0111010: q = 4'b1000;
		10'b010_0111011: q = 4'b1000;
		10'b010_0111100: q = 4'b1000;
		10'b010_0111101: q = 4'b1000;
		10'b010_0111110: q = 4'b1000;
		10'b010_0111111: q = 4'b1000;
		10'b010_1000000: q = 4'b0001;
		10'b010_1000001: q = 4'b0001;
		10'b010_1000010: q = 4'b0001;
		10'b010_1000011: q = 4'b0001;
		10'b010_1000100: q = 4'b0001;
		10'b010_1000101: q = 4'b0001;
		10'b010_1000110: q = 4'b0001;
		10'b010_1000111: q = 4'b0001;
		10'b010_1001000: q = 4'b0001;
		10'b010_1001001: q = 4'b0001;
		10'b010_1001010: q = 4'b0001;
		10'b010_1001011: q = 4'b0001;
		10'b010_1001100: q = 4'b0001;
		10'b010_1001101: q = 4'b0001;
		10'b010_1001110: q = 4'b0001;
		10'b010_1001111: q = 4'b0001;
		10'b010_1010000: q = 4'b0001;
		10'b010_1010001: q = 4'b0001;
		10'b010_1010010: q = 4'b0001;
		10'b010_1010011: q = 4'b0001;
		10'b010_1010100: q = 4'b0001;
		10'b010_1010101: q = 4'b0001;
		10'b010_1010110: q = 4'b0001;
		10'b010_1010111: q = 4'b0001;
		10'b010_1011000: q = 4'b0001;
		10'b010_1011001: q = 4'b0001;
		10'b010_1011010: q = 4'b0001;
		10'b010_1011011: q = 4'b0001;
		10'b010_1011100: q = 4'b0001;
		10'b010_1011101: q = 4'b0001;
		10'b010_1011110: q = 4'b0001;
		10'b010_1011111: q = 4'b0001;
		10'b010_1100000: q = 4'b0001;
		10'b010_1100001: q = 4'b0001;
		10'b010_1100010: q = 4'b0001;
		10'b010_1100011: q = 4'b0001;
		10'b010_1100100: q = 4'b0001;
		10'b010_1100101: q = 4'b0001;
		10'b010_1100110: q = 4'b0001;
		10'b010_1100111: q = 4'b0001;
		10'b010_1101000: q = 4'b0001;
		10'b010_1101001: q = 4'b0001;
		10'b010_1101010: q = 4'b0001;
		10'b010_1101011: q = 4'b0001;
		10'b010_1101100: q = 4'b0001;
		10'b010_1101101: q = 4'b0001;
		10'b010_1101110: q = 4'b0001;
		10'b010_1101111: q = 4'b0001;
		10'b010_1110000: q = 4'b0010;
		10'b010_1110001: q = 4'b0010;
		10'b010_1110010: q = 4'b0010;
		10'b010_1110011: q = 4'b0010;
		10'b010_1110100: q = 4'b0010;
		10'b010_1110101: q = 4'b0010;
		10'b010_1110110: q = 4'b0010;
		10'b010_1110111: q = 4'b0010;
		10'b010_1111000: q = 4'b0010;
		10'b010_1111001: q = 4'b0010;
		10'b010_1111010: q = 4'b0000;
		10'b010_1111011: q = 4'b0000;
		10'b010_1111100: q = 4'b0000;
		10'b010_1111101: q = 4'b0000;
		10'b010_1111110: q = 4'b0000;
		10'b010_1111111: q = 4'b0000;
		10'b011_0000000: q = 4'b0000;
		10'b011_0000001: q = 4'b0000;
		10'b011_0000010: q = 4'b0000;
		10'b011_0000011: q = 4'b0000;
		10'b011_0000100: q = 4'b0100;
		10'b011_0000101: q = 4'b0100;
		10'b011_0000110: q = 4'b0100;
		10'b011_0000111: q = 4'b0100;
		10'b011_0001000: q = 4'b0100;
		10'b011_0001001: q = 4'b0100;
		10'b011_0001010: q = 4'b0100;
		10'b011_0001011: q = 4'b0100;
		10'b011_0001100: q = 4'b0100;
		10'b011_0001101: q = 4'b0100;
		10'b011_0001110: q = 4'b0100;
		10'b011_0001111: q = 4'b0100;
		10'b011_0010000: q = 4'b1000;
		10'b011_0010001: q = 4'b1000;
		10'b011_0010010: q = 4'b1000;
		10'b011_0010011: q = 4'b1000;
		10'b011_0010100: q = 4'b1000;
		10'b011_0010101: q = 4'b1000;
		10'b011_0010110: q = 4'b1000;
		10'b011_0010111: q = 4'b1000;
		10'b011_0011000: q = 4'b1000;
		10'b011_0011001: q = 4'b1000;
		10'b011_0011010: q = 4'b1000;
		10'b011_0011011: q = 4'b1000;
		10'b011_0011100: q = 4'b1000;
		10'b011_0011101: q = 4'b1000;
		10'b011_0011110: q = 4'b1000;
		10'b011_0011111: q = 4'b1000;
		10'b011_0100000: q = 4'b1000;
		10'b011_0100001: q = 4'b1000;
		10'b011_0100010: q = 4'b1000;
		10'b011_0100011: q = 4'b1000;
		10'b011_0100100: q = 4'b1000;
		10'b011_0100101: q = 4'b1000;
		10'b011_0100110: q = 4'b1000;
		10'b011_0100111: q = 4'b1000;
		10'b011_0101000: q = 4'b1000;
		10'b011_0101001: q = 4'b1000;
		10'b011_0101010: q = 4'b1000;
		10'b011_0101011: q = 4'b1000;
		10'b011_0101100: q = 4'b1000;
		10'b011_0101101: q = 4'b1000;
		10'b011_0101110: q = 4'b1000;
		10'b011_0101111: q = 4'b1000;
		10'b011_0110000: q = 4'b1000;
		10'b011_0110001: q = 4'b1000;
		10'b011_0110010: q = 4'b1000;
		10'b011_0110011: q = 4'b1000;
		10'b011_0110100: q = 4'b1000;
		10'b011_0110101: q = 4'b1000;
		10'b011_0110110: q = 4'b1000;
		10'b011_0110111: q = 4'b1000;
		10'b011_0111000: q = 4'b1000;
		10'b011_0111001: q = 4'b1000;
		10'b011_0111010: q = 4'b1000;
		10'b011_0111011: q = 4'b1000;
		10'b011_0111100: q = 4'b1000;
		10'b011_0111101: q = 4'b1000;
		10'b011_0111110: q = 4'b1000;
		10'b011_0111111: q = 4'b1000;
		10'b011_1000000: q = 4'b0001;
		10'b011_1000001: q = 4'b0001;
		10'b011_1000010: q = 4'b0001;
		10'b011_1000011: q = 4'b0001;
		10'b011_1000100: q = 4'b0001;
		10'b011_1000101: q = 4'b0001;
		10'b011_1000110: q = 4'b0001;
		10'b011_1000111: q = 4'b0001;
		10'b011_1001000: q = 4'b0001;
		10'b011_1001001: q = 4'b0001;
		10'b011_1001010: q = 4'b0001;
		10'b011_1001011: q = 4'b0001;
		10'b011_1001100: q = 4'b0001;
		10'b011_1001101: q = 4'b0001;
		10'b011_1001110: q = 4'b0001;
		10'b011_1001111: q = 4'b0001;
		10'b011_1010000: q = 4'b0001;
		10'b011_1010001: q = 4'b0001;
		10'b011_1010010: q = 4'b0001;
		10'b011_1010011: q = 4'b0001;
		10'b011_1010100: q = 4'b0001;
		10'b011_1010101: q = 4'b0001;
		10'b011_1010110: q = 4'b0001;
		10'b011_1010111: q = 4'b0001;
		10'b011_1011000: q = 4'b0001;
		10'b011_1011001: q = 4'b0001;
		10'b011_1011010: q = 4'b0001;
		10'b011_1011011: q = 4'b0001;
		10'b011_1011100: q = 4'b0001;
		10'b011_1011101: q = 4'b0001;
		10'b011_1011110: q = 4'b0001;
		10'b011_1011111: q = 4'b0001;
		10'b011_1100000: q = 4'b0001;
		10'b011_1100001: q = 4'b0001;
		10'b011_1100010: q = 4'b0001;
		10'b011_1100011: q = 4'b0001;
		10'b011_1100100: q = 4'b0001;
		10'b011_1100101: q = 4'b0001;
		10'b011_1100110: q = 4'b0001;
		10'b011_1100111: q = 4'b0001;
		10'b011_1101000: q = 4'b0001;
		10'b011_1101001: q = 4'b0001;
		10'b011_1101010: q = 4'b0001;
		10'b011_1101011: q = 4'b0001;
		10'b011_1101100: q = 4'b0001;
		10'b011_1101101: q = 4'b0001;
		10'b011_1101110: q = 4'b0010;
		10'b011_1101111: q = 4'b0010;
		10'b011_1110000: q = 4'b0010;
		10'b011_1110001: q = 4'b0010;
		10'b011_1110010: q = 4'b0010;
		10'b011_1110011: q = 4'b0010;
		10'b011_1110100: q = 4'b0010;
		10'b011_1110101: q = 4'b0010;
		10'b011_1110110: q = 4'b0010;
		10'b011_1110111: q = 4'b0010;
		10'b011_1111000: q = 4'b0010;
		10'b011_1111001: q = 4'b0010;
		10'b011_1111010: q = 4'b0000;
		10'b011_1111011: q = 4'b0000;
		10'b011_1111100: q = 4'b0000;
		10'b011_1111101: q = 4'b0000;
		10'b011_1111110: q = 4'b0000;
		10'b011_1111111: q = 4'b0000;
		10'b100_0000000: q = 4'b0000;
		10'b100_0000001: q = 4'b0000;
		10'b100_0000010: q = 4'b0000;
		10'b100_0000011: q = 4'b0000;
		10'b100_0000100: q = 4'b0000;
		10'b100_0000101: q = 4'b0000;
		10'b100_0000110: q = 4'b0100;
		10'b100_0000111: q = 4'b0100;
		10'b100_0001000: q = 4'b0100;
		10'b100_0001001: q = 4'b0100;
		10'b100_0001010: q = 4'b0100;
		10'b100_0001011: q = 4'b0100;
		10'b100_0001100: q = 4'b0100;
		10'b100_0001101: q = 4'b0100;
		10'b100_0001110: q = 4'b0100;
		10'b100_0001111: q = 4'b0100;
		10'b100_0010000: q = 4'b0100;
		10'b100_0010001: q = 4'b0100;
		10'b100_0010010: q = 4'b1000;
		10'b100_0010011: q = 4'b1000;
		10'b100_0010100: q = 4'b1000;
		10'b100_0010101: q = 4'b1000;
		10'b100_0010110: q = 4'b1000;
		10'b100_0010111: q = 4'b1000;
		10'b100_0011000: q = 4'b1000;
		10'b100_0011001: q = 4'b1000;
		10'b100_0011010: q = 4'b1000;
		10'b100_0011011: q = 4'b1000;
		10'b100_0011100: q = 4'b1000;
		10'b100_0011101: q = 4'b1000;
		10'b100_0011110: q = 4'b1000;
		10'b100_0011111: q = 4'b1000;
		10'b100_0100000: q = 4'b1000;
		10'b100_0100001: q = 4'b1000;
		10'b100_0100010: q = 4'b1000;
		10'b100_0100011: q = 4'b1000;
		10'b100_0100100: q = 4'b1000;
		10'b100_0100101: q = 4'b1000;
		10'b100_0100110: q = 4'b1000;
		10'b100_0100111: q = 4'b1000;
		10'b100_0101000: q = 4'b1000;
		10'b100_0101001: q = 4'b1000;
		10'b100_0101010: q = 4'b1000;
		10'b100_0101011: q = 4'b1000;
		10'b100_0101100: q = 4'b1000;
		10'b100_0101101: q = 4'b1000;
		10'b100_0101110: q = 4'b1000;
		10'b100_0101111: q = 4'b1000;
		10'b100_0110000: q = 4'b1000;
		10'b100_0110001: q = 4'b1000;
		10'b100_0110010: q = 4'b1000;
		10'b100_0110011: q = 4'b1000;
		10'b100_0110100: q = 4'b1000;
		10'b100_0110101: q = 4'b1000;
		10'b100_0110110: q = 4'b1000;
		10'b100_0110111: q = 4'b1000;
		10'b100_0111000: q = 4'b1000;
		10'b100_0111001: q = 4'b1000;
		10'b100_0111010: q = 4'b1000;
		10'b100_0111011: q = 4'b1000;
		10'b100_0111100: q = 4'b1000;
		10'b100_0111101: q = 4'b1000;
		10'b100_0111110: q = 4'b1000;
		10'b100_0111111: q = 4'b1000;
		10'b100_1000000: q = 4'b0001;
		10'b100_1000001: q = 4'b0001;
		10'b100_1000010: q = 4'b0001;
		10'b100_1000011: q = 4'b0001;
		10'b100_1000100: q = 4'b0001;
		10'b100_1000101: q = 4'b0001;
		10'b100_1000110: q = 4'b0001;
		10'b100_1000111: q = 4'b0001;
		10'b100_1001000: q = 4'b0001;
		10'b100_1001001: q = 4'b0001;
		10'b100_1001010: q = 4'b0001;
		10'b100_1001011: q = 4'b0001;
		10'b100_1001100: q = 4'b0001;
		10'b100_1001101: q = 4'b0001;
		10'b100_1001110: q = 4'b0001;
		10'b100_1001111: q = 4'b0001;
		10'b100_1010000: q = 4'b0001;
		10'b100_1010001: q = 4'b0001;
		10'b100_1010010: q = 4'b0001;
		10'b100_1010011: q = 4'b0001;
		10'b100_1010100: q = 4'b0001;
		10'b100_1010101: q = 4'b0001;
		10'b100_1010110: q = 4'b0001;
		10'b100_1010111: q = 4'b0001;
		10'b100_1011000: q = 4'b0001;
		10'b100_1011001: q = 4'b0001;
		10'b100_1011010: q = 4'b0001;
		10'b100_1011011: q = 4'b0001;
		10'b100_1011100: q = 4'b0001;
		10'b100_1011101: q = 4'b0001;
		10'b100_1011110: q = 4'b0001;
		10'b100_1011111: q = 4'b0001;
		10'b100_1100000: q = 4'b0001;
		10'b100_1100001: q = 4'b0001;
		10'b100_1100010: q = 4'b0001;
		10'b100_1100011: q = 4'b0001;
		10'b100_1100100: q = 4'b0001;
		10'b100_1100101: q = 4'b0001;
		10'b100_1100110: q = 4'b0001;
		10'b100_1100111: q = 4'b0001;
		10'b100_1101000: q = 4'b0001;
		10'b100_1101001: q = 4'b0001;
		10'b100_1101010: q = 4'b0001;
		10'b100_1101011: q = 4'b0001;
		10'b100_1101100: q = 4'b0010;
		10'b100_1101101: q = 4'b0010;
		10'b100_1101110: q = 4'b0010;
		10'b100_1101111: q = 4'b0010;
		10'b100_1110000: q = 4'b0010;
		10'b100_1110001: q = 4'b0010;
		10'b100_1110010: q = 4'b0010;
		10'b100_1110011: q = 4'b0010;
		10'b100_1110100: q = 4'b0010;
		10'b100_1110101: q = 4'b0010;
		10'b100_1110110: q = 4'b0010;
		10'b100_1110111: q = 4'b0010;
		10'b100_1111000: q = 4'b0000;
		10'b100_1111001: q = 4'b0000;
		10'b100_1111010: q = 4'b0000;
		10'b100_1111011: q = 4'b0000;
		10'b100_1111100: q = 4'b0000;
		10'b100_1111101: q = 4'b0000;
		10'b100_1111110: q = 4'b0000;
		10'b100_1111111: q = 4'b0000;
		10'b101_0000000: q = 4'b0000;
		10'b101_0000001: q = 4'b0000;
		10'b101_0000010: q = 4'b0000;
		10'b101_0000011: q = 4'b0000;
		10'b101_0000100: q = 4'b0000;
		10'b101_0000101: q = 4'b0000;
		10'b101_0000110: q = 4'b0100;
		10'b101_0000111: q = 4'b0100;
		10'b101_0001000: q = 4'b0100;
		10'b101_0001001: q = 4'b0100;
		10'b101_0001010: q = 4'b0100;
		10'b101_0001011: q = 4'b0100;
		10'b101_0001100: q = 4'b0100;
		10'b101_0001101: q = 4'b0100;
		10'b101_0001110: q = 4'b0100;
		10'b101_0001111: q = 4'b0100;
		10'b101_0010000: q = 4'b0100;
		10'b101_0010001: q = 4'b0100;
		10'b101_0010010: q = 4'b0100;
		10'b101_0010011: q = 4'b0100;
		10'b101_0010100: q = 4'b1000;
		10'b101_0010101: q = 4'b1000;
		10'b101_0010110: q = 4'b1000;
		10'b101_0010111: q = 4'b1000;
		10'b101_0011000: q = 4'b1000;
		10'b101_0011001: q = 4'b1000;
		10'b101_0011010: q = 4'b1000;
		10'b101_0011011: q = 4'b1000;
		10'b101_0011100: q = 4'b1000;
		10'b101_0011101: q = 4'b1000;
		10'b101_0011110: q = 4'b1000;
		10'b101_0011111: q = 4'b1000;
		10'b101_0100000: q = 4'b1000;
		10'b101_0100001: q = 4'b1000;
		10'b101_0100010: q = 4'b1000;
		10'b101_0100011: q = 4'b1000;
		10'b101_0100100: q = 4'b1000;
		10'b101_0100101: q = 4'b1000;
		10'b101_0100110: q = 4'b1000;
		10'b101_0100111: q = 4'b1000;
		10'b101_0101000: q = 4'b1000;
		10'b101_0101001: q = 4'b1000;
		10'b101_0101010: q = 4'b1000;
		10'b101_0101011: q = 4'b1000;
		10'b101_0101100: q = 4'b1000;
		10'b101_0101101: q = 4'b1000;
		10'b101_0101110: q = 4'b1000;
		10'b101_0101111: q = 4'b1000;
		10'b101_0110000: q = 4'b1000;
		10'b101_0110001: q = 4'b1000;
		10'b101_0110010: q = 4'b1000;
		10'b101_0110011: q = 4'b1000;
		10'b101_0110100: q = 4'b1000;
		10'b101_0110101: q = 4'b1000;
		10'b101_0110110: q = 4'b1000;
		10'b101_0110111: q = 4'b1000;
		10'b101_0111000: q = 4'b1000;
		10'b101_0111001: q = 4'b1000;
		10'b101_0111010: q = 4'b1000;
		10'b101_0111011: q = 4'b1000;
		10'b101_0111100: q = 4'b1000;
		10'b101_0111101: q = 4'b1000;
		10'b101_0111110: q = 4'b1000;
		10'b101_0111111: q = 4'b1000;
		10'b101_1000000: q = 4'b0001;
		10'b101_1000001: q = 4'b0001;
		10'b101_1000010: q = 4'b0001;
		10'b101_1000011: q = 4'b0001;
		10'b101_1000100: q = 4'b0001;
		10'b101_1000101: q = 4'b0001;
		10'b101_1000110: q = 4'b0001;
		10'b101_1000111: q = 4'b0001;
		10'b101_1001000: q = 4'b0001;
		10'b101_1001001: q = 4'b0001;
		10'b101_1001010: q = 4'b0001;
		10'b101_1001011: q = 4'b0001;
		10'b101_1001100: q = 4'b0001;
		10'b101_1001101: q = 4'b0001;
		10'b101_1001110: q = 4'b0001;
		10'b101_1001111: q = 4'b0001;
		10'b101_1010000: q = 4'b0001;
		10'b101_1010001: q = 4'b0001;
		10'b101_1010010: q = 4'b0001;
		10'b101_1010011: q = 4'b0001;
		10'b101_1010100: q = 4'b0001;
		10'b101_1010101: q = 4'b0001;
		10'b101_1010110: q = 4'b0001;
		10'b101_1010111: q = 4'b0001;
		10'b101_1011000: q = 4'b0001;
		10'b101_1011001: q = 4'b0001;
		10'b101_1011010: q = 4'b0001;
		10'b101_1011011: q = 4'b0001;
		10'b101_1011100: q = 4'b0001;
		10'b101_1011101: q = 4'b0001;
		10'b101_1011110: q = 4'b0001;
		10'b101_1011111: q = 4'b0001;
		10'b101_1100000: q = 4'b0001;
		10'b101_1100001: q = 4'b0001;
		10'b101_1100010: q = 4'b0001;
		10'b101_1100011: q = 4'b0001;
		10'b101_1100100: q = 4'b0001;
		10'b101_1100101: q = 4'b0001;
		10'b101_1100110: q = 4'b0001;
		10'b101_1100111: q = 4'b0001;
		10'b101_1101000: q = 4'b0001;
		10'b101_1101001: q = 4'b0001;
		10'b101_1101010: q = 4'b0001;
		10'b101_1101011: q = 4'b0001;
		10'b101_1101100: q = 4'b0010;
		10'b101_1101101: q = 4'b0010;
		10'b101_1101110: q = 4'b0010;
		10'b101_1101111: q = 4'b0010;
		10'b101_1110000: q = 4'b0010;
		10'b101_1110001: q = 4'b0010;
		10'b101_1110010: q = 4'b0010;
		10'b101_1110011: q = 4'b0010;
		10'b101_1110100: q = 4'b0010;
		10'b101_1110101: q = 4'b0010;
		10'b101_1110110: q = 4'b0010;
		10'b101_1110111: q = 4'b0010;
		10'b101_1111000: q = 4'b0000;
		10'b101_1111001: q = 4'b0000;
		10'b101_1111010: q = 4'b0000;
		10'b101_1111011: q = 4'b0000;
		10'b101_1111100: q = 4'b0000;
		10'b101_1111101: q = 4'b0000;
		10'b101_1111110: q = 4'b0000;
		10'b101_1111111: q = 4'b0000;
		10'b110_0000000: q = 4'b0000;
		10'b110_0000001: q = 4'b0000;
		10'b110_0000010: q = 4'b0000;
		10'b110_0000011: q = 4'b0000;
		10'b110_0000100: q = 4'b0000;
		10'b110_0000101: q = 4'b0000;
		10'b110_0000110: q = 4'b0000;
		10'b110_0000111: q = 4'b0000;
		10'b110_0001000: q = 4'b0100;
		10'b110_0001001: q = 4'b0100;
		10'b110_0001010: q = 4'b0100;
		10'b110_0001011: q = 4'b0100;
		10'b110_0001100: q = 4'b0100;
		10'b110_0001101: q = 4'b0100;
		10'b110_0001110: q = 4'b0100;
		10'b110_0001111: q = 4'b0100;
		10'b110_0010000: q = 4'b0100;
		10'b110_0010001: q = 4'b0100;
		10'b110_0010010: q = 4'b0100;
		10'b110_0010011: q = 4'b0100;
		10'b110_0010100: q = 4'b1000;
		10'b110_0010101: q = 4'b1000;
		10'b110_0010110: q = 4'b1000;
		10'b110_0010111: q = 4'b1000;
		10'b110_0011000: q = 4'b1000;
		10'b110_0011001: q = 4'b1000;
		10'b110_0011010: q = 4'b1000;
		10'b110_0011011: q = 4'b1000;
		10'b110_0011100: q = 4'b1000;
		10'b110_0011101: q = 4'b1000;
		10'b110_0011110: q = 4'b1000;
		10'b110_0011111: q = 4'b1000;
		10'b110_0100000: q = 4'b1000;
		10'b110_0100001: q = 4'b1000;
		10'b110_0100010: q = 4'b1000;
		10'b110_0100011: q = 4'b1000;
		10'b110_0100100: q = 4'b1000;
		10'b110_0100101: q = 4'b1000;
		10'b110_0100110: q = 4'b1000;
		10'b110_0100111: q = 4'b1000;
		10'b110_0101000: q = 4'b1000;
		10'b110_0101001: q = 4'b1000;
		10'b110_0101010: q = 4'b1000;
		10'b110_0101011: q = 4'b1000;
		10'b110_0101100: q = 4'b1000;
		10'b110_0101101: q = 4'b1000;
		10'b110_0101110: q = 4'b1000;
		10'b110_0101111: q = 4'b1000;
		10'b110_0110000: q = 4'b1000;
		10'b110_0110001: q = 4'b1000;
		10'b110_0110010: q = 4'b1000;
		10'b110_0110011: q = 4'b1000;
		10'b110_0110100: q = 4'b1000;
		10'b110_0110101: q = 4'b1000;
		10'b110_0110110: q = 4'b1000;
		10'b110_0110111: q = 4'b1000;
		10'b110_0111000: q = 4'b1000;
		10'b110_0111001: q = 4'b1000;
		10'b110_0111010: q = 4'b1000;
		10'b110_0111011: q = 4'b1000;
		10'b110_0111100: q = 4'b1000;
		10'b110_0111101: q = 4'b1000;
		10'b110_0111110: q = 4'b1000;
		10'b110_0111111: q = 4'b1000;
		10'b110_1000000: q = 4'b0001;
		10'b110_1000001: q = 4'b0001;
		10'b110_1000010: q = 4'b0001;
		10'b110_1000011: q = 4'b0001;
		10'b110_1000100: q = 4'b0001;
		10'b110_1000101: q = 4'b0001;
		10'b110_1000110: q = 4'b0001;
		10'b110_1000111: q = 4'b0001;
		10'b110_1001000: q = 4'b0001;
		10'b110_1001001: q = 4'b0001;
		10'b110_1001010: q = 4'b0001;
		10'b110_1001011: q = 4'b0001;
		10'b110_1001100: q = 4'b0001;
		10'b110_1001101: q = 4'b0001;
		10'b110_1001110: q = 4'b0001;
		10'b110_1001111: q = 4'b0001;
		10'b110_1010000: q = 4'b0001;
		10'b110_1010001: q = 4'b0001;
		10'b110_1010010: q = 4'b0001;
		10'b110_1010011: q = 4'b0001;
		10'b110_1010100: q = 4'b0001;
		10'b110_1010101: q = 4'b0001;
		10'b110_1010110: q = 4'b0001;
		10'b110_1010111: q = 4'b0001;
		10'b110_1011000: q = 4'b0001;
		10'b110_1011001: q = 4'b0001;
		10'b110_1011010: q = 4'b0001;
		10'b110_1011011: q = 4'b0001;
		10'b110_1011100: q = 4'b0001;
		10'b110_1011101: q = 4'b0001;
		10'b110_1011110: q = 4'b0001;
		10'b110_1011111: q = 4'b0001;
		10'b110_1100000: q = 4'b0001;
		10'b110_1100001: q = 4'b0001;
		10'b110_1100010: q = 4'b0001;
		10'b110_1100011: q = 4'b0001;
		10'b110_1100100: q = 4'b0001;
		10'b110_1100101: q = 4'b0001;
		10'b110_1100110: q = 4'b0001;
		10'b110_1100111: q = 4'b0001;
		10'b110_1101000: q = 4'b0001;
		10'b110_1101001: q = 4'b0001;
		10'b110_1101010: q = 4'b0010;
		10'b110_1101011: q = 4'b0010;
		10'b110_1101100: q = 4'b0010;
		10'b110_1101101: q = 4'b0010;
		10'b110_1101110: q = 4'b0010;
		10'b110_1101111: q = 4'b0010;
		10'b110_1110000: q = 4'b0010;
		10'b110_1110001: q = 4'b0010;
		10'b110_1110010: q = 4'b0010;
		10'b110_1110011: q = 4'b0010;
		10'b110_1110100: q = 4'b0010;
		10'b110_1110101: q = 4'b0010;
		10'b110_1110110: q = 4'b0010;
		10'b110_1110111: q = 4'b0010;
		10'b110_1111000: q = 4'b0000;
		10'b110_1111001: q = 4'b0000;
		10'b110_1111010: q = 4'b0000;
		10'b110_1111011: q = 4'b0000;
		10'b110_1111100: q = 4'b0000;
		10'b110_1111101: q = 4'b0000;
		10'b110_1111110: q = 4'b0000;
		10'b110_1111111: q = 4'b0000;
		10'b111_0000000: q = 4'b0000;
		10'b111_0000001: q = 4'b0000;
		10'b111_0000010: q = 4'b0000;
		10'b111_0000011: q = 4'b0000;
		10'b111_0000100: q = 4'b0000;
		10'b111_0000101: q = 4'b0000;
		10'b111_0000110: q = 4'b0000;
		10'b111_0000111: q = 4'b0000;
		10'b111_0001000: q = 4'b0100;
		10'b111_0001001: q = 4'b0100;
		10'b111_0001010: q = 4'b0100;
		10'b111_0001011: q = 4'b0100;
		10'b111_0001100: q = 4'b0100;
		10'b111_0001101: q = 4'b0100;
		10'b111_0001110: q = 4'b0100;
		10'b111_0001111: q = 4'b0100;
		10'b111_0010000: q = 4'b0100;
		10'b111_0010001: q = 4'b0100;
		10'b111_0010010: q = 4'b0100;
		10'b111_0010011: q = 4'b0100;
		10'b111_0010100: q = 4'b0100;
		10'b111_0010101: q = 4'b0100;
		10'b111_0010110: q = 4'b0100;
		10'b111_0010111: q = 4'b0100;
		10'b111_0011000: q = 4'b1000;
		10'b111_0011001: q = 4'b1000;
		10'b111_0011010: q = 4'b1000;
		10'b111_0011011: q = 4'b1000;
		10'b111_0011100: q = 4'b1000;
		10'b111_0011101: q = 4'b1000;
		10'b111_0011110: q = 4'b1000;
		10'b111_0011111: q = 4'b1000;
		10'b111_0100000: q = 4'b1000;
		10'b111_0100001: q = 4'b1000;
		10'b111_0100010: q = 4'b1000;
		10'b111_0100011: q = 4'b1000;
		10'b111_0100100: q = 4'b1000;
		10'b111_0100101: q = 4'b1000;
		10'b111_0100110: q = 4'b1000;
		10'b111_0100111: q = 4'b1000;
		10'b111_0101000: q = 4'b1000;
		10'b111_0101001: q = 4'b1000;
		10'b111_0101010: q = 4'b1000;
		10'b111_0101011: q = 4'b1000;
		10'b111_0101100: q = 4'b1000;
		10'b111_0101101: q = 4'b1000;
		10'b111_0101110: q = 4'b1000;
		10'b111_0101111: q = 4'b1000;
		10'b111_0110000: q = 4'b1000;
		10'b111_0110001: q = 4'b1000;
		10'b111_0110010: q = 4'b1000;
		10'b111_0110011: q = 4'b1000;
		10'b111_0110100: q = 4'b1000;
		10'b111_0110101: q = 4'b1000;
		10'b111_0110110: q = 4'b1000;
		10'b111_0110111: q = 4'b1000;
		10'b111_0111000: q = 4'b1000;
		10'b111_0111001: q = 4'b1000;
		10'b111_0111010: q = 4'b1000;
		10'b111_0111011: q = 4'b1000;
		10'b111_0111100: q = 4'b1000;
		10'b111_0111101: q = 4'b1000;
		10'b111_0111110: q = 4'b1000;
		10'b111_0111111: q = 4'b1000;
		10'b111_1000000: q = 4'b0001;
		10'b111_1000001: q = 4'b0001;
		10'b111_1000010: q = 4'b0001;
		10'b111_1000011: q = 4'b0001;
		10'b111_1000100: q = 4'b0001;
		10'b111_1000101: q = 4'b0001;
		10'b111_1000110: q = 4'b0001;
		10'b111_1000111: q = 4'b0001;
		10'b111_1001000: q = 4'b0001;
		10'b111_1001001: q = 4'b0001;
		10'b111_1001010: q = 4'b0001;
		10'b111_1001011: q = 4'b0001;
		10'b111_1001100: q = 4'b0001;
		10'b111_1001101: q = 4'b0001;
		10'b111_1001110: q = 4'b0001;
		10'b111_1001111: q = 4'b0001;
		10'b111_1010000: q = 4'b0001;
		10'b111_1010001: q = 4'b0001;
		10'b111_1010010: q = 4'b0001;
		10'b111_1010011: q = 4'b0001;
		10'b111_1010100: q = 4'b0001;
		10'b111_1010101: q = 4'b0001;
		10'b111_1010110: q = 4'b0001;
		10'b111_1010111: q = 4'b0001;
		10'b111_1011000: q = 4'b0001;
		10'b111_1011001: q = 4'b0001;
		10'b111_1011010: q = 4'b0001;
		10'b111_1011011: q = 4'b0001;
		10'b111_1011100: q = 4'b0001;
		10'b111_1011101: q = 4'b0001;
		10'b111_1011110: q = 4'b0001;
		10'b111_1011111: q = 4'b0001;
		10'b111_1100000: q = 4'b0001;
		10'b111_1100001: q = 4'b0001;
		10'b111_1100010: q = 4'b0001;
		10'b111_1100011: q = 4'b0001;
		10'b111_1100100: q = 4'b0001;
		10'b111_1100101: q = 4'b0001;
		10'b111_1100110: q = 4'b0001;
		10'b111_1100111: q = 4'b0001;
		10'b111_1101000: q = 4'b0010;
		10'b111_1101001: q = 4'b0010;
		10'b111_1101010: q = 4'b0010;
		10'b111_1101011: q = 4'b0010;
		10'b111_1101100: q = 4'b0010;
		10'b111_1101101: q = 4'b0010;
		10'b111_1101110: q = 4'b0010;
		10'b111_1101111: q = 4'b0010;
		10'b111_1110000: q = 4'b0010;
		10'b111_1110001: q = 4'b0010;
		10'b111_1110010: q = 4'b0010;
		10'b111_1110011: q = 4'b0010;
		10'b111_1110100: q = 4'b0010;
		10'b111_1110101: q = 4'b0010;
		10'b111_1110110: q = 4'b0010;
		10'b111_1110111: q = 4'b0010;
		10'b111_1111000: q = 4'b0000;
		10'b111_1111001: q = 4'b0000;
		10'b111_1111010: q = 4'b0000;
		10'b111_1111011: q = 4'b0000;
		10'b111_1111100: q = 4'b0000;
		10'b111_1111101: q = 4'b0000;
		10'b111_1111110: q = 4'b0000;
		10'b111_1111111: q = 4'b0000;
	endcase

endmodule
///////////////////////////////////////////
// galoismult_forward.sv
//
// Written: ryan.swann@okstate.edu, james.stine@okstate.edu, David_Harris@hmc.edu
// Created: 20 February 2024
//
// Purpose: Galois field operations for mix columns operation
//
// A component of the CORE-V-WALLY configurable RISC-V project.
// https://github.com/openhwgroup/cvw
// 
// Copyright (C) 2021-24 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

module galoismult_forward (
   input  logic [7:0] in,
   output logic [7:0] out);

   logic [7:0] leftshift;

   assign leftshift = {in[6:0], 1'b0};
   assign out = in[7] ? (leftshift ^ 8'b00011011) : leftshift;

endmodule

module gm2 (gm2_In, gm2_Out); 
   
   input logic [7:0]  gm2_In;
   output logic [7:0] gm2_Out;
   
   // Set output to Galois Mult 2
   assign gm2_Out = {gm2_In[6:0], 1'b0} ^ (8'h1b & {8{gm2_In[7]}});
   
endmodule 
///////////////////////////////////////////
//
// Written: James Stine
// Modified: 8/1/2018
//
// Purpose: Bipartite Lookup
// 
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// MIT LICENSE
// Permission is hereby granted, free of charge, to any person obtaining a copy of this 
// software and associated documentation files (the "Software"), to deal in the Software 
// without restriction, including without limitation the rights to use, copy, modify, merge, 
// publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons 
// to whom the Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in all copies or 
//   substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, 
//   INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR 
//   PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS 
//   BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, 
//   TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE 
//   OR OTHER DEALINGS IN THE SOFTWARE.
////////////////////////////////////////////////////////////////////////////////////////////////

module sbtm_a3 (input  logic [7:0] a,
		output logic [5:0] y);
   
   always_comb
     case(a)
       8'b01000000: y = 6'b100110;
       8'b01000001: y = 6'b100001;
       8'b01000010: y = 6'b011100;
       8'b01000011: y = 6'b010111;
       8'b01000100: y = 6'b010010;
       8'b01000101: y = 6'b001100;
       8'b01000110: y = 6'b000111;
       8'b01000111: y = 6'b000010;
       8'b01001000: y = 6'b100000;
       8'b01001001: y = 6'b011100;
       8'b01001010: y = 6'b011000;
       8'b01001011: y = 6'b010011;
       8'b01001100: y = 6'b001111;
       8'b01001101: y = 6'b001010;
       8'b01001110: y = 6'b000110;
       8'b01001111: y = 6'b000010;
       8'b01010000: y = 6'b011100;
       8'b01010001: y = 6'b011000;
       8'b01010010: y = 6'b010100;
       8'b01010011: y = 6'b010000;
       8'b01010100: y = 6'b001101;
       8'b01010101: y = 6'b001001;
       8'b01010110: y = 6'b000101;
       8'b01010111: y = 6'b000001;
       8'b01011000: y = 6'b011000;
       8'b01011001: y = 6'b010101;
       8'b01011010: y = 6'b010010;
       8'b01011011: y = 6'b001110;
       8'b01011100: y = 6'b001011;
       8'b01011101: y = 6'b001000;
       8'b01011110: y = 6'b000100;
       8'b01011111: y = 6'b000001;
       8'b01100000: y = 6'b010101;
       8'b01100001: y = 6'b010010;
       8'b01100010: y = 6'b001111;
       8'b01100011: y = 6'b001101;
       8'b01100100: y = 6'b001010;
       8'b01100101: y = 6'b000111;
       8'b01100110: y = 6'b000100;
       8'b01100111: y = 6'b000001;
       8'b01101000: y = 6'b010011;
       8'b01101001: y = 6'b010000;
       8'b01101010: y = 6'b001110;
       8'b01101011: y = 6'b001011;
       8'b01101100: y = 6'b001001;
       8'b01101101: y = 6'b000110;
       8'b01101110: y = 6'b000011;
       8'b01101111: y = 6'b000001;
       8'b01110000: y = 6'b010001;
       8'b01110001: y = 6'b001111;
       8'b01110010: y = 6'b001100;
       8'b01110011: y = 6'b001010;
       8'b01110100: y = 6'b001000;
       8'b01110101: y = 6'b000101;
       8'b01110110: y = 6'b000011;
       8'b01110111: y = 6'b000001;
       8'b01111000: y = 6'b001111;
       8'b01111001: y = 6'b001101;
       8'b01111010: y = 6'b001011;
       8'b01111011: y = 6'b001001;
       8'b01111100: y = 6'b000111;
       8'b01111101: y = 6'b000101;
       8'b01111110: y = 6'b000011;
       8'b01111111: y = 6'b000001;       
       8'b10000000: y = 6'b001110;
       8'b10000001: y = 6'b001100;
       8'b10000010: y = 6'b001010;
       8'b10000011: y = 6'b001000;
       8'b10000100: y = 6'b000110;
       8'b10000101: y = 6'b000100;
       8'b10000110: y = 6'b000010;
       8'b10000111: y = 6'b000000;
       8'b10001000: y = 6'b001101;
       8'b10001001: y = 6'b001011;
       8'b10001010: y = 6'b001001;
       8'b10001011: y = 6'b000111;
       8'b10001100: y = 6'b000110;
       8'b10001101: y = 6'b000100;
       8'b10001110: y = 6'b000010;
       8'b10001111: y = 6'b000000;
       8'b10010000: y = 6'b001100;
       8'b10010001: y = 6'b001010;
       8'b10010010: y = 6'b001000;
       8'b10010011: y = 6'b000111;
       8'b10010100: y = 6'b000101;
       8'b10010101: y = 6'b000100;
       8'b10010110: y = 6'b000010;
       8'b10010111: y = 6'b000000;
       8'b10011000: y = 6'b001011;
       8'b10011001: y = 6'b001001;
       8'b10011010: y = 6'b001000;
       8'b10011011: y = 6'b000110;
       8'b10011100: y = 6'b000101;
       8'b10011101: y = 6'b000011;
       8'b10011110: y = 6'b000010;
       8'b10011111: y = 6'b000000;
       8'b10100000: y = 6'b001010;
       8'b10100001: y = 6'b001000;
       8'b10100010: y = 6'b000111;
       8'b10100011: y = 6'b000110;
       8'b10100100: y = 6'b000100;
       8'b10100101: y = 6'b000011;
       8'b10100110: y = 6'b000010;
       8'b10100111: y = 6'b000000;
       8'b10101000: y = 6'b001001;
       8'b10101001: y = 6'b001000;
       8'b10101010: y = 6'b000111;
       8'b10101011: y = 6'b000101;
       8'b10101100: y = 6'b000100;
       8'b10101101: y = 6'b000011;
       8'b10101110: y = 6'b000001;
       8'b10101111: y = 6'b000000;
       8'b10110000: y = 6'b001000;
       8'b10110001: y = 6'b000111;
       8'b10110010: y = 6'b000110;
       8'b10110011: y = 6'b000101;
       8'b10110100: y = 6'b000100;
       8'b10110101: y = 6'b000010;
       8'b10110110: y = 6'b000001;
       8'b10110111: y = 6'b000000;
       8'b10111000: y = 6'b001000;
       8'b10111001: y = 6'b000111;
       8'b10111010: y = 6'b000110;
       8'b10111011: y = 6'b000101;
       8'b10111100: y = 6'b000011;
       8'b10111101: y = 6'b000010;
       8'b10111110: y = 6'b000001;
       8'b10111111: y = 6'b000000;
       8'b11000000: y = 6'b000111;
       8'b11000001: y = 6'b000110;
       8'b11000010: y = 6'b000101;
       8'b11000011: y = 6'b000100;
       8'b11000100: y = 6'b000011;
       8'b11000101: y = 6'b000010;
       8'b11000110: y = 6'b000001;
       8'b11000111: y = 6'b000000;
       8'b11001000: y = 6'b000111;
       8'b11001001: y = 6'b000110;
       8'b11001010: y = 6'b000101;
       8'b11001011: y = 6'b000100;
       8'b11001100: y = 6'b000011;
       8'b11001101: y = 6'b000010;
       8'b11001110: y = 6'b000001;
       8'b11001111: y = 6'b000000;
       8'b11010000: y = 6'b000111;
       8'b11010001: y = 6'b000110;
       8'b11010010: y = 6'b000101;
       8'b11010011: y = 6'b000100;
       8'b11010100: y = 6'b000011;
       8'b11010101: y = 6'b000010;
       8'b11010110: y = 6'b000001;
       8'b11010111: y = 6'b000000;
       8'b11011000: y = 6'b000110;
       8'b11011001: y = 6'b000101;
       8'b11011010: y = 6'b000100;
       8'b11011011: y = 6'b000011;
       8'b11011100: y = 6'b000011;
       8'b11011101: y = 6'b000010;
       8'b11011110: y = 6'b000001;
       8'b11011111: y = 6'b000000;
       8'b11100000: y = 6'b000110;
       8'b11100001: y = 6'b000101;
       8'b11100010: y = 6'b000100;
       8'b11100011: y = 6'b000011;
       8'b11100100: y = 6'b000010;
       8'b11100101: y = 6'b000010;
       8'b11100110: y = 6'b000001;
       8'b11100111: y = 6'b000000;
       8'b11101000: y = 6'b000101;
       8'b11101001: y = 6'b000101;
       8'b11101010: y = 6'b000100;
       8'b11101011: y = 6'b000011;
       8'b11101100: y = 6'b000010;
       8'b11101101: y = 6'b000001;
       8'b11101110: y = 6'b000001;
       8'b11101111: y = 6'b000000;
       8'b11110000: y = 6'b000101;
       8'b11110001: y = 6'b000100;
       8'b11110010: y = 6'b000100;
       8'b11110011: y = 6'b000011;
       8'b11110100: y = 6'b000010;
       8'b11110101: y = 6'b000001;
       8'b11110110: y = 6'b000001;
       8'b11110111: y = 6'b000000;
       8'b11111000: y = 6'b000101;
       8'b11111001: y = 6'b000100;
       8'b11111010: y = 6'b000011;
       8'b11111011: y = 6'b000011;
       8'b11111100: y = 6'b000010;
       8'b11111101: y = 6'b000001;
       8'b11111110: y = 6'b000001;
       8'b11111111: y = 6'b000000;
       default: y = 6'bxxxxxx;
     endcase // case (a)
    
endmodule // sbtm_a0

// Brent-Kung Carry-save Prefix Adder

module bk128 (cout, sum, a, b, cin);
   
   input [127:0] a, b;
   input 	 cin;
   
   output [127:0] sum;
   output 	  cout;

   wire [128:0]   p,g,t;
   wire [127:0]   c;

   // pre-computation
   assign p={a^b,1'b0};
   assign g={a&b, cin};
   assign t[1]=p[1];
   assign t[2]=p[2];
   assign t[3]=p[3]^g[2];
   assign t[4]=p[4];
   assign t[5]=p[5]^g[4];
   assign t[6]=p[6];
   assign t[7]=p[7]^g[6];
   assign t[8]=p[8];
   assign t[9]=p[9]^g[8];
   assign t[10]=p[10];
   assign t[11]=p[11]^g[10];
   assign t[12]=p[12];
   assign t[13]=p[13]^g[12];
   assign t[14]=p[14];
   assign t[15]=p[15]^g[14];
   assign t[16]=p[16];
   assign t[17]=p[17]^g[16];
   assign t[18]=p[18];
   assign t[19]=p[19]^g[18];
   assign t[20]=p[20];
   assign t[21]=p[21]^g[20];
   assign t[22]=p[22];
   assign t[23]=p[23]^g[22];
   assign t[24]=p[24];
   assign t[25]=p[25]^g[24];
   assign t[26]=p[26];
   assign t[27]=p[27]^g[26];
   assign t[28]=p[28];
   assign t[29]=p[29]^g[28];
   assign t[30]=p[30];
   assign t[31]=p[31]^g[30];
   assign t[32]=p[32];
   assign t[33]=p[33]^g[32];
   assign t[34]=p[34];
   assign t[35]=p[35]^g[34];
   assign t[36]=p[36];
   assign t[37]=p[37]^g[36];
   assign t[38]=p[38];
   assign t[39]=p[39]^g[38];
   assign t[40]=p[40];
   assign t[41]=p[41]^g[40];
   assign t[42]=p[42];
   assign t[43]=p[43]^g[42];
   assign t[44]=p[44];
   assign t[45]=p[45]^g[44];
   assign t[46]=p[46];
   assign t[47]=p[47]^g[46];
   assign t[48]=p[48];
   assign t[49]=p[49]^g[48];
   assign t[50]=p[50];
   assign t[51]=p[51]^g[50];
   assign t[52]=p[52];
   assign t[53]=p[53]^g[52];
   assign t[54]=p[54];
   assign t[55]=p[55]^g[54];
   assign t[56]=p[56];
   assign t[57]=p[57]^g[56];
   assign t[58]=p[58];
   assign t[59]=p[59]^g[58];
   assign t[60]=p[60];
   assign t[61]=p[61]^g[60];
   assign t[62]=p[62];
   assign t[63]=p[63]^g[62];
   assign t[64]=p[64];
   assign t[65]=p[65]^g[64];
   assign t[66]=p[66];
   assign t[67]=p[67]^g[66];
   assign t[68]=p[68];
   assign t[69]=p[69]^g[68];
   assign t[70]=p[70];
   assign t[71]=p[71]^g[70];
   assign t[72]=p[72];
   assign t[73]=p[73]^g[72];
   assign t[74]=p[74];
   assign t[75]=p[75]^g[74];
   assign t[76]=p[76];
   assign t[77]=p[77]^g[76];
   assign t[78]=p[78];
   assign t[79]=p[79]^g[78];
   assign t[80]=p[80];
   assign t[81]=p[81]^g[80];
   assign t[82]=p[82];
   assign t[83]=p[83]^g[82];
   assign t[84]=p[84];
   assign t[85]=p[85]^g[84];
   assign t[86]=p[86];
   assign t[87]=p[87]^g[86];
   assign t[88]=p[88];
   assign t[89]=p[89]^g[88];
   assign t[90]=p[90];
   assign t[91]=p[91]^g[90];
   assign t[92]=p[92];
   assign t[93]=p[93]^g[92];
   assign t[94]=p[94];
   assign t[95]=p[95]^g[94];
   assign t[96]=p[96];
   assign t[97]=p[97]^g[96];
   assign t[98]=p[98];
   assign t[99]=p[99]^g[98];
   assign t[100]=p[100];
   assign t[101]=p[101]^g[100];
   assign t[102]=p[102];
   assign t[103]=p[103]^g[102];
   assign t[104]=p[104];
   assign t[105]=p[105]^g[104];
   assign t[106]=p[106];
   assign t[107]=p[107]^g[106];
   assign t[108]=p[108];
   assign t[109]=p[109]^g[108];
   assign t[110]=p[110];
   assign t[111]=p[111]^g[110];
   assign t[112]=p[112];
   assign t[113]=p[113]^g[112];
   assign t[114]=p[114];
   assign t[115]=p[115]^g[114];
   assign t[116]=p[116];
   assign t[117]=p[117]^g[116];
   assign t[118]=p[118];
   assign t[119]=p[119]^g[118];
   assign t[120]=p[120];
   assign t[121]=p[121]^g[120];
   assign t[122]=p[122];
   assign t[123]=p[123]^g[122];
   assign t[124]=p[124];
   assign t[125]=p[125]^g[124];
   assign t[126]=p[126];
   assign t[127]=p[127]^g[126];
   assign t[128]=p[128];

   // prefix tree
   brent_kung_cs128 prefix_tree(c, p[127:0], g[127:0]);

   // post-computation
   assign sum=p[128:1]^c;
   assign cout=g[128]|(p[128]&c[127]);

endmodule

module brent_kung_cs128 (c, p, g);
   
   input [127:0] p;
   input [127:0] g;
   output [128:1] c;


   // parallel-prefix, Brent-Kung

   // Stage 1: Generates G/P pairs that span 1 bits
   grey b_1_0 (G_1_0, {g[1],g[0]}, p[1]);
   black b_3_2 (G_3_2, P_3_2, {g[3],g[2]}, {p[3],p[2]});
   black b_5_4 (G_5_4, P_5_4, {g[5],g[4]}, {p[5],p[4]});
   black b_7_6 (G_7_6, P_7_6, {g[7],g[6]}, {p[7],p[6]});
   black b_9_8 (G_9_8, P_9_8, {g[9],g[8]}, {p[9],p[8]});
   black b_11_10 (G_11_10, P_11_10, {g[11],g[10]}, {p[11],p[10]});
   black b_13_12 (G_13_12, P_13_12, {g[13],g[12]}, {p[13],p[12]});
   black b_15_14 (G_15_14, P_15_14, {g[15],g[14]}, {p[15],p[14]});

   black b_17_16 (G_17_16, P_17_16, {g[17],g[16]}, {p[17],p[16]});
   black b_19_18 (G_19_18, P_19_18, {g[19],g[18]}, {p[19],p[18]});
   black b_21_20 (G_21_20, P_21_20, {g[21],g[20]}, {p[21],p[20]});
   black b_23_22 (G_23_22, P_23_22, {g[23],g[22]}, {p[23],p[22]});
   black b_25_24 (G_25_24, P_25_24, {g[25],g[24]}, {p[25],p[24]});
   black b_27_26 (G_27_26, P_27_26, {g[27],g[26]}, {p[27],p[26]});
   black b_29_28 (G_29_28, P_29_28, {g[29],g[28]}, {p[29],p[28]});
   black b_31_30 (G_31_30, P_31_30, {g[31],g[30]}, {p[31],p[30]});

   black b_33_32 (G_33_32, P_33_32, {g[33],g[32]}, {p[33],p[32]});
   black b_35_34 (G_35_34, P_35_34, {g[35],g[34]}, {p[35],p[34]});
   black b_37_36 (G_37_36, P_37_36, {g[37],g[36]}, {p[37],p[36]});
   black b_39_38 (G_39_38, P_39_38, {g[39],g[38]}, {p[39],p[38]});
   black b_41_40 (G_41_40, P_41_40, {g[41],g[40]}, {p[41],p[40]});
   black b_43_42 (G_43_42, P_43_42, {g[43],g[42]}, {p[43],p[42]});
   black b_45_44 (G_45_44, P_45_44, {g[45],g[44]}, {p[45],p[44]});
   black b_47_46 (G_47_46, P_47_46, {g[47],g[46]}, {p[47],p[46]});

   black b_49_48 (G_49_48, P_49_48, {g[49],g[48]}, {p[49],p[48]});
   black b_51_50 (G_51_50, P_51_50, {g[51],g[50]}, {p[51],p[50]});
   black b_53_52 (G_53_52, P_53_52, {g[53],g[52]}, {p[53],p[52]});
   black b_55_54 (G_55_54, P_55_54, {g[55],g[54]}, {p[55],p[54]});
   black b_57_56 (G_57_56, P_57_56, {g[57],g[56]}, {p[57],p[56]});
   black b_59_58 (G_59_58, P_59_58, {g[59],g[58]}, {p[59],p[58]});
   black b_61_60 (G_61_60, P_61_60, {g[61],g[60]}, {p[61],p[60]});
   black b_63_62 (G_63_62, P_63_62, {g[63],g[62]}, {p[63],p[62]});

   black b_65_64 (G_65_64, P_65_64, {g[65],g[64]}, {p[65],p[64]});
   black b_67_66 (G_67_66, P_67_66, {g[67],g[66]}, {p[67],p[66]});
   black b_69_68 (G_69_68, P_69_68, {g[69],g[68]}, {p[69],p[68]});
   black b_71_70 (G_71_70, P_71_70, {g[71],g[70]}, {p[71],p[70]});
   black b_73_72 (G_73_72, P_73_72, {g[73],g[72]}, {p[73],p[72]});
   black b_75_74 (G_75_74, P_75_74, {g[75],g[74]}, {p[75],p[74]});
   black b_77_76 (G_77_76, P_77_76, {g[77],g[76]}, {p[77],p[76]});
   black b_79_78 (G_79_78, P_79_78, {g[79],g[78]}, {p[79],p[78]});

   black b_81_80 (G_81_80, P_81_80, {g[81],g[80]}, {p[81],p[80]});
   black b_83_82 (G_83_82, P_83_82, {g[83],g[82]}, {p[83],p[82]});
   black b_85_84 (G_85_84, P_85_84, {g[85],g[84]}, {p[85],p[84]});
   black b_87_86 (G_87_86, P_87_86, {g[87],g[86]}, {p[87],p[86]});
   black b_89_88 (G_89_88, P_89_88, {g[89],g[88]}, {p[89],p[88]});
   black b_91_90 (G_91_90, P_91_90, {g[91],g[90]}, {p[91],p[90]});
   black b_93_92 (G_93_92, P_93_92, {g[93],g[92]}, {p[93],p[92]});
   black b_95_94 (G_95_94, P_95_94, {g[95],g[94]}, {p[95],p[94]});

   black b_97_96 (G_97_96, P_97_96, {g[97],g[96]}, {p[97],p[96]});
   black b_99_98 (G_99_98, P_99_98, {g[99],g[98]}, {p[99],p[98]});
   black b_101_100 (G_101_100, P_101_100, {g[101],g[100]}, {p[101],p[100]});
   black b_103_102 (G_103_102, P_103_102, {g[103],g[102]}, {p[103],p[102]});
   black b_105_104 (G_105_104, P_105_104, {g[105],g[104]}, {p[105],p[104]});
   black b_107_106 (G_107_106, P_107_106, {g[107],g[106]}, {p[107],p[106]});
   black b_109_108 (G_109_108, P_109_108, {g[109],g[108]}, {p[109],p[108]});
   black b_111_110 (G_111_110, P_111_110, {g[111],g[110]}, {p[111],p[110]});

   black b_113_112 (G_113_112, P_113_112, {g[113],g[112]}, {p[113],p[112]});
   black b_115_114 (G_115_114, P_115_114, {g[115],g[114]}, {p[115],p[114]});
   black b_117_116 (G_117_116, P_117_116, {g[117],g[116]}, {p[117],p[116]});
   black b_119_118 (G_119_118, P_119_118, {g[119],g[118]}, {p[119],p[118]});
   black b_121_120 (G_121_120, P_121_120, {g[121],g[120]}, {p[121],p[120]});
   black b_123_122 (G_123_122, P_123_122, {g[123],g[122]}, {p[123],p[122]});
   black b_125_124 (G_125_124, P_125_124, {g[125],g[124]}, {p[125],p[124]});
   black b_127_126 (G_127_126, P_127_126, {g[127],g[126]}, {p[127],p[126]});


   // Stage 2: Generates G/P pairs that span 2 bits
   grey g_3_0 (G_3_0, {G_3_2,G_1_0}, P_3_2);
   black b_7_4 (G_7_4, P_7_4, {G_7_6,G_5_4}, {P_7_6,P_5_4});
   black b_11_8 (G_11_8, P_11_8, {G_11_10,G_9_8}, {P_11_10,P_9_8});
   black b_15_12 (G_15_12, P_15_12, {G_15_14,G_13_12}, {P_15_14,P_13_12});
   black b_19_16 (G_19_16, P_19_16, {G_19_18,G_17_16}, {P_19_18,P_17_16});
   black b_23_20 (G_23_20, P_23_20, {G_23_22,G_21_20}, {P_23_22,P_21_20});
   black b_27_24 (G_27_24, P_27_24, {G_27_26,G_25_24}, {P_27_26,P_25_24});
   black b_31_28 (G_31_28, P_31_28, {G_31_30,G_29_28}, {P_31_30,P_29_28});

   black b_35_32 (G_35_32, P_35_32, {G_35_34,G_33_32}, {P_35_34,P_33_32});
   black b_39_36 (G_39_36, P_39_36, {G_39_38,G_37_36}, {P_39_38,P_37_36});
   black b_43_40 (G_43_40, P_43_40, {G_43_42,G_41_40}, {P_43_42,P_41_40});
   black b_47_44 (G_47_44, P_47_44, {G_47_46,G_45_44}, {P_47_46,P_45_44});
   black b_51_48 (G_51_48, P_51_48, {G_51_50,G_49_48}, {P_51_50,P_49_48});
   black b_55_52 (G_55_52, P_55_52, {G_55_54,G_53_52}, {P_55_54,P_53_52});
   black b_59_56 (G_59_56, P_59_56, {G_59_58,G_57_56}, {P_59_58,P_57_56});
   black b_63_60 (G_63_60, P_63_60, {G_63_62,G_61_60}, {P_63_62,P_61_60});

   black b_67_64 (G_67_64, P_67_64, {G_67_66,G_65_64}, {P_67_66,P_65_64});
   black b_71_68 (G_71_68, P_71_68, {G_71_70,G_69_68}, {P_71_70,P_69_68});
   black b_75_72 (G_75_72, P_75_72, {G_75_74,G_73_72}, {P_75_74,P_73_72});
   black b_79_76 (G_79_76, P_79_76, {G_79_78,G_77_76}, {P_79_78,P_77_76});
   black b_83_80 (G_83_80, P_83_80, {G_83_82,G_81_80}, {P_83_82,P_81_80});
   black b_87_84 (G_87_84, P_87_84, {G_87_86,G_85_84}, {P_87_86,P_85_84});
   black b_91_88 (G_91_88, P_91_88, {G_91_90,G_89_88}, {P_91_90,P_89_88});
   black b_95_92 (G_95_92, P_95_92, {G_95_94,G_93_92}, {P_95_94,P_93_92});

   black b_99_96 (G_99_96, P_99_96, {G_99_98,G_97_96}, {P_99_98,P_97_96});
   black b_103_100 (G_103_100, P_103_100, {G_103_102,G_101_100}, {P_103_102,P_101_100});
   black b_107_104 (G_107_104, P_107_104, {G_107_106,G_105_104}, {P_107_106,P_105_104});
   black b_111_108 (G_111_108, P_111_108, {G_111_110,G_109_108}, {P_111_110,P_109_108});
   black b_115_112 (G_115_112, P_115_112, {G_115_114,G_113_112}, {P_115_114,P_113_112});
   black b_119_116 (G_119_116, P_119_116, {G_119_118,G_117_116}, {P_119_118,P_117_116});
   black b_123_120 (G_123_120, P_123_120, {G_123_122,G_121_120}, {P_123_122,P_121_120});
   black b_127_124 (G_127_124, P_127_124, {G_127_126,G_125_124}, {P_127_126,P_125_124});


   // Stage 3: Generates G/P pairs that span 4 bits
   grey g_7_0 (G_7_0, {G_7_4,G_3_0}, P_7_4);
   black b_15_8 (G_15_8, P_15_8, {G_15_12,G_11_8}, {P_15_12,P_11_8});
   black b_23_16 (G_23_16, P_23_16, {G_23_20,G_19_16}, {P_23_20,P_19_16});
   black b_31_24 (G_31_24, P_31_24, {G_31_28,G_27_24}, {P_31_28,P_27_24});
   black b_39_32 (G_39_32, P_39_32, {G_39_36,G_35_32}, {P_39_36,P_35_32});
   black b_47_40 (G_47_40, P_47_40, {G_47_44,G_43_40}, {P_47_44,P_43_40});
   black b_55_48 (G_55_48, P_55_48, {G_55_52,G_51_48}, {P_55_52,P_51_48});
   black b_63_56 (G_63_56, P_63_56, {G_63_60,G_59_56}, {P_63_60,P_59_56});

   black b_71_64 (G_71_64, P_71_64, {G_71_68,G_67_64}, {P_71_68,P_67_64});
   black b_79_72 (G_79_72, P_79_72, {G_79_76,G_75_72}, {P_79_76,P_75_72});
   black b_87_80 (G_87_80, P_87_80, {G_87_84,G_83_80}, {P_87_84,P_83_80});
   black b_95_88 (G_95_88, P_95_88, {G_95_92,G_91_88}, {P_95_92,P_91_88});
   black b_103_96 (G_103_96, P_103_96, {G_103_100,G_99_96}, {P_103_100,P_99_96});
   black b_111_104 (G_111_104, P_111_104, {G_111_108,G_107_104}, {P_111_108,P_107_104});
   black b_119_112 (G_119_112, P_119_112, {G_119_116,G_115_112}, {P_119_116,P_115_112});
   black b_127_120 (G_127_120, P_127_120, {G_127_124,G_123_120}, {P_127_124,P_123_120});


   // Stage 4: Generates G/P pairs that span 8 bits
   grey g_15_0 (G_15_0, {G_15_8,G_7_0}, P_15_8);
   black b_31_16 (G_31_16, P_31_16, {G_31_24,G_23_16}, {P_31_24,P_23_16});
   black b_47_32 (G_47_32, P_47_32, {G_47_40,G_39_32}, {P_47_40,P_39_32});
   black b_63_48 (G_63_48, P_63_48, {G_63_56,G_55_48}, {P_63_56,P_55_48});
   black b_79_64 (G_79_64, P_79_64, {G_79_72,G_71_64}, {P_79_72,P_71_64});
   black b_95_80 (G_95_80, P_95_80, {G_95_88,G_87_80}, {P_95_88,P_87_80});
   black b_111_96 (G_111_96, P_111_96, {G_111_104,G_103_96}, {P_111_104,P_103_96});
   black b_127_112 (G_127_112, P_127_112, {G_127_120,G_119_112}, {P_127_120,P_119_112});


   // Stage 5: Generates G/P pairs that span 16 bits
   grey g_31_0 (G_31_0, {G_31_16,G_15_0}, P_31_16);
   black b_63_32 (G_63_32, P_63_32, {G_63_48,G_47_32}, {P_63_48,P_47_32});
   black b_95_64 (G_95_64, P_95_64, {G_95_80,G_79_64}, {P_95_80,P_79_64});
   black b_127_96 (G_127_96, P_127_96, {G_127_112,G_111_96}, {P_127_112,P_111_96});

   // Stage 6: Generates G/P pairs that span 32 bits
   grey g_63_0 (G_63_0, {G_63_32,G_31_0}, P_63_32);
   black b_127_64 (G_127_64, P_127_64, {G_127_96,G_95_64}, {P_127_96,P_95_64});

   // Stage 7: Generates G/P pairs that span 64 bits
   grey g_127_0 (G_127_0, {G_127_64,G_63_0}, P_127_64);

   // Stage 8: Generates G/P pairs that span 32 bits
   grey g_95_0 (G_95_0, {G_95_64,G_63_0}, P_95_64);

   // Stage 9: Generates G/P pairs that span 16 bits
   grey g_47_0 (G_47_0, {G_47_32,G_31_0}, P_47_32);
   grey g_79_0 (G_79_0, {G_79_64,G_63_0}, P_79_64);
   grey g_111_0 (G_111_0, {G_111_96,G_95_0}, P_111_96);

   // Stage 10: Generates G/P pairs that span 8 bits
   grey g_23_0 (G_23_0, {G_23_16,G_15_0}, P_23_16);
   grey g_39_0 (G_39_0, {G_39_32,G_31_0}, P_39_32);
   grey g_55_0 (G_55_0, {G_55_48,G_47_0}, P_55_48);
   grey g_71_0 (G_71_0, {G_71_64,G_63_0}, P_71_64);
   grey g_87_0 (G_87_0, {G_87_80,G_79_0}, P_87_80);
   grey g_103_0 (G_103_0, {G_103_96,G_95_0}, P_103_96);
   grey g_119_0 (G_119_0, {G_119_112,G_111_0}, P_119_112);

   // Stage 11: Generates G/P pairs that span 4 bits
   grey g_11_0 (G_11_0, {G_11_8,G_7_0}, P_11_8);
   grey g_19_0 (G_19_0, {G_19_16,G_15_0}, P_19_16);
   grey g_27_0 (G_27_0, {G_27_24,G_23_0}, P_27_24);
   grey g_35_0 (G_35_0, {G_35_32,G_31_0}, P_35_32);
   grey g_43_0 (G_43_0, {G_43_40,G_39_0}, P_43_40);
   grey g_51_0 (G_51_0, {G_51_48,G_47_0}, P_51_48);
   grey g_59_0 (G_59_0, {G_59_56,G_55_0}, P_59_56);
   grey g_67_0 (G_67_0, {G_67_64,G_63_0}, P_67_64);
   grey g_75_0 (G_75_0, {G_75_72,G_71_0}, P_75_72);
   grey g_83_0 (G_83_0, {G_83_80,G_79_0}, P_83_80);
   grey g_91_0 (G_91_0, {G_91_88,G_87_0}, P_91_88);
   grey g_99_0 (G_99_0, {G_99_96,G_95_0}, P_99_96);
   grey g_107_0 (G_107_0, {G_107_104,G_103_0}, P_107_104);
   grey g_115_0 (G_115_0, {G_115_112,G_111_0}, P_115_112);
   grey g_123_0 (G_123_0, {G_123_120,G_119_0}, P_123_120);

   // Stage 12: Generates G/P pairs that span 2 bits
   grey g_5_0 (G_5_0, {G_5_4,G_3_0}, P_5_4);
   grey g_9_0 (G_9_0, {G_9_8,G_7_0}, P_9_8);
   grey g_13_0 (G_13_0, {G_13_12,G_11_0}, P_13_12);
   grey g_17_0 (G_17_0, {G_17_16,G_15_0}, P_17_16);
   grey g_21_0 (G_21_0, {G_21_20,G_19_0}, P_21_20);
   grey g_25_0 (G_25_0, {G_25_24,G_23_0}, P_25_24);
   grey g_29_0 (G_29_0, {G_29_28,G_27_0}, P_29_28);
   grey g_33_0 (G_33_0, {G_33_32,G_31_0}, P_33_32);
   grey g_37_0 (G_37_0, {G_37_36,G_35_0}, P_37_36);
   grey g_41_0 (G_41_0, {G_41_40,G_39_0}, P_41_40);
   grey g_45_0 (G_45_0, {G_45_44,G_43_0}, P_45_44);
   grey g_49_0 (G_49_0, {G_49_48,G_47_0}, P_49_48);
   grey g_53_0 (G_53_0, {G_53_52,G_51_0}, P_53_52);
   grey g_57_0 (G_57_0, {G_57_56,G_55_0}, P_57_56);
   grey g_61_0 (G_61_0, {G_61_60,G_59_0}, P_61_60);
   grey g_65_0 (G_65_0, {G_65_64,G_63_0}, P_65_64);
   grey g_69_0 (G_69_0, {G_69_68,G_67_0}, P_69_68);
   grey g_73_0 (G_73_0, {G_73_72,G_71_0}, P_73_72);
   grey g_77_0 (G_77_0, {G_77_76,G_75_0}, P_77_76);
   grey g_81_0 (G_81_0, {G_81_80,G_79_0}, P_81_80);
   grey g_85_0 (G_85_0, {G_85_84,G_83_0}, P_85_84);
   grey g_89_0 (G_89_0, {G_89_88,G_87_0}, P_89_88);
   grey g_93_0 (G_93_0, {G_93_92,G_91_0}, P_93_92);
   grey g_97_0 (G_97_0, {G_97_96,G_95_0}, P_97_96);
   grey g_101_0 (G_101_0, {G_101_100,G_99_0}, P_101_100);
   grey g_105_0 (G_105_0, {G_105_104,G_103_0}, P_105_104);
   grey g_109_0 (G_109_0, {G_109_108,G_107_0}, P_109_108);
   grey g_113_0 (G_113_0, {G_113_112,G_111_0}, P_113_112);
   grey g_117_0 (G_117_0, {G_117_116,G_115_0}, P_117_116);
   grey g_121_0 (G_121_0, {G_121_120,G_119_0}, P_121_120);
   grey g_125_0 (G_125_0, {G_125_124,G_123_0}, P_125_124);

   // Last grey cell stage 
   grey g_2_0 (G_2_0, {g[2],G_1_0}, p[2]);
   grey g_4_0 (G_4_0, {g[4],G_3_0}, p[4]);
   grey g_6_0 (G_6_0, {g[6],G_5_0}, p[6]);
   grey g_8_0 (G_8_0, {g[8],G_7_0}, p[8]);
   grey g_10_0 (G_10_0, {g[10],G_9_0}, p[10]);
   grey g_12_0 (G_12_0, {g[12],G_11_0}, p[12]);
   grey g_14_0 (G_14_0, {g[14],G_13_0}, p[14]);
   grey g_16_0 (G_16_0, {g[16],G_15_0}, p[16]);
   grey g_18_0 (G_18_0, {g[18],G_17_0}, p[18]);
   grey g_20_0 (G_20_0, {g[20],G_19_0}, p[20]);
   grey g_22_0 (G_22_0, {g[22],G_21_0}, p[22]);
   grey g_24_0 (G_24_0, {g[24],G_23_0}, p[24]);
   grey g_26_0 (G_26_0, {g[26],G_25_0}, p[26]);
   grey g_28_0 (G_28_0, {g[28],G_27_0}, p[28]);
   grey g_30_0 (G_30_0, {g[30],G_29_0}, p[30]);
   grey g_32_0 (G_32_0, {g[32],G_31_0}, p[32]);
   grey g_34_0 (G_34_0, {g[34],G_33_0}, p[34]);
   grey g_36_0 (G_36_0, {g[36],G_35_0}, p[36]);
   grey g_38_0 (G_38_0, {g[38],G_37_0}, p[38]);
   grey g_40_0 (G_40_0, {g[40],G_39_0}, p[40]);
   grey g_42_0 (G_42_0, {g[42],G_41_0}, p[42]);
   grey g_44_0 (G_44_0, {g[44],G_43_0}, p[44]);
   grey g_46_0 (G_46_0, {g[46],G_45_0}, p[46]);
   grey g_48_0 (G_48_0, {g[48],G_47_0}, p[48]);
   grey g_50_0 (G_50_0, {g[50],G_49_0}, p[50]);
   grey g_52_0 (G_52_0, {g[52],G_51_0}, p[52]);
   grey g_54_0 (G_54_0, {g[54],G_53_0}, p[54]);
   grey g_56_0 (G_56_0, {g[56],G_55_0}, p[56]);
   grey g_58_0 (G_58_0, {g[58],G_57_0}, p[58]);
   grey g_60_0 (G_60_0, {g[60],G_59_0}, p[60]);
   grey g_62_0 (G_62_0, {g[62],G_61_0}, p[62]);
   grey g_64_0 (G_64_0, {g[64],G_63_0}, p[64]);
   grey g_66_0 (G_66_0, {g[66],G_65_0}, p[66]);
   grey g_68_0 (G_68_0, {g[68],G_67_0}, p[68]);
   grey g_70_0 (G_70_0, {g[70],G_69_0}, p[70]);
   grey g_72_0 (G_72_0, {g[72],G_71_0}, p[72]);
   grey g_74_0 (G_74_0, {g[74],G_73_0}, p[74]);
   grey g_76_0 (G_76_0, {g[76],G_75_0}, p[76]);
   grey g_78_0 (G_78_0, {g[78],G_77_0}, p[78]);
   grey g_80_0 (G_80_0, {g[80],G_79_0}, p[80]);
   grey g_82_0 (G_82_0, {g[82],G_81_0}, p[82]);
   grey g_84_0 (G_84_0, {g[84],G_83_0}, p[84]);
   grey g_86_0 (G_86_0, {g[86],G_85_0}, p[86]);
   grey g_88_0 (G_88_0, {g[88],G_87_0}, p[88]);
   grey g_90_0 (G_90_0, {g[90],G_89_0}, p[90]);
   grey g_92_0 (G_92_0, {g[92],G_91_0}, p[92]);
   grey g_94_0 (G_94_0, {g[94],G_93_0}, p[94]);
   grey g_96_0 (G_96_0, {g[96],G_95_0}, p[96]);
   grey g_98_0 (G_98_0, {g[98],G_97_0}, p[98]);
   grey g_100_0 (G_100_0, {g[100],G_99_0}, p[100]);
   grey g_102_0 (G_102_0, {g[102],G_101_0}, p[102]);
   grey g_104_0 (G_104_0, {g[104],G_103_0}, p[104]);
   grey g_106_0 (G_106_0, {g[106],G_105_0}, p[106]);
   grey g_108_0 (G_108_0, {g[108],G_107_0}, p[108]);
   grey g_110_0 (G_110_0, {g[110],G_109_0}, p[110]);
   grey g_112_0 (G_112_0, {g[112],G_111_0}, p[112]);
   grey g_114_0 (G_114_0, {g[114],G_113_0}, p[114]);
   grey g_116_0 (G_116_0, {g[116],G_115_0}, p[116]);
   grey g_118_0 (G_118_0, {g[118],G_117_0}, p[118]);
   grey g_120_0 (G_120_0, {g[120],G_119_0}, p[120]);
   grey g_122_0 (G_122_0, {g[122],G_121_0}, p[122]);
   grey g_124_0 (G_124_0, {g[124],G_123_0}, p[124]);
   grey g_126_0 (G_126_0, {g[126],G_125_0}, p[126]);

   // Final Stage: Apply c_k+1=G_k_0
   assign c[1]=g[0];
   assign c[2]=G_1_0;
   assign c[3]=G_2_0;
   assign c[4]=G_3_0;
   assign c[5]=G_4_0;
   assign c[6]=G_5_0;
   assign c[7]=G_6_0;
   assign c[8]=G_7_0;
   assign c[9]=G_8_0;

   assign c[10]=G_9_0;
   assign c[11]=G_10_0;
   assign c[12]=G_11_0;
   assign c[13]=G_12_0;
   assign c[14]=G_13_0;
   assign c[15]=G_14_0;
   assign c[16]=G_15_0;
   assign c[17]=G_16_0;

   assign c[18]=G_17_0;
   assign c[19]=G_18_0;
   assign c[20]=G_19_0;
   assign c[21]=G_20_0;
   assign c[22]=G_21_0;
   assign c[23]=G_22_0;
   assign c[24]=G_23_0;
   assign c[25]=G_24_0;

   assign c[26]=G_25_0;
   assign c[27]=G_26_0;
   assign c[28]=G_27_0;
   assign c[29]=G_28_0;
   assign c[30]=G_29_0;
   assign c[31]=G_30_0;
   assign c[32]=G_31_0;
   assign c[33]=G_32_0;

   assign c[34]=G_33_0;
   assign c[35]=G_34_0;
   assign c[36]=G_35_0;
   assign c[37]=G_36_0;
   assign c[38]=G_37_0;
   assign c[39]=G_38_0;
   assign c[40]=G_39_0;
   assign c[41]=G_40_0;

   assign c[42]=G_41_0;
   assign c[43]=G_42_0;
   assign c[44]=G_43_0;
   assign c[45]=G_44_0;
   assign c[46]=G_45_0;
   assign c[47]=G_46_0;
   assign c[48]=G_47_0;
   assign c[49]=G_48_0;

   assign c[50]=G_49_0;
   assign c[51]=G_50_0;
   assign c[52]=G_51_0;
   assign c[53]=G_52_0;
   assign c[54]=G_53_0;
   assign c[55]=G_54_0;
   assign c[56]=G_55_0;
   assign c[57]=G_56_0;

   assign c[58]=G_57_0;
   assign c[59]=G_58_0;
   assign c[60]=G_59_0;
   assign c[61]=G_60_0;
   assign c[62]=G_61_0;
   assign c[63]=G_62_0;
   assign c[64]=G_63_0;
   assign c[65]=G_64_0;

   assign c[66]=G_65_0;
   assign c[67]=G_66_0;
   assign c[68]=G_67_0;
   assign c[69]=G_68_0;
   assign c[70]=G_69_0;
   assign c[71]=G_70_0;
   assign c[72]=G_71_0;
   assign c[73]=G_72_0;

   assign c[74]=G_73_0;
   assign c[75]=G_74_0;
   assign c[76]=G_75_0;
   assign c[77]=G_76_0;
   assign c[78]=G_77_0;
   assign c[79]=G_78_0;
   assign c[80]=G_79_0;
   assign c[81]=G_80_0;

   assign c[82]=G_81_0;
   assign c[83]=G_82_0;
   assign c[84]=G_83_0;
   assign c[85]=G_84_0;
   assign c[86]=G_85_0;
   assign c[87]=G_86_0;
   assign c[88]=G_87_0;
   assign c[89]=G_88_0;

   assign c[90]=G_89_0;
   assign c[91]=G_90_0;
   assign c[92]=G_91_0;
   assign c[93]=G_92_0;
   assign c[94]=G_93_0;
   assign c[95]=G_94_0;
   assign c[96]=G_95_0;
   assign c[97]=G_96_0;

   assign c[98]=G_97_0;
   assign c[99]=G_98_0;
   assign c[100]=G_99_0;
   assign c[101]=G_100_0;
   assign c[102]=G_101_0;
   assign c[103]=G_102_0;
   assign c[104]=G_103_0;
   assign c[105]=G_104_0;

   assign c[106]=G_105_0;
   assign c[107]=G_106_0;
   assign c[108]=G_107_0;
   assign c[109]=G_108_0;
   assign c[110]=G_109_0;
   assign c[111]=G_110_0;
   assign c[112]=G_111_0;
   assign c[113]=G_112_0;

   assign c[114]=G_113_0;
   assign c[115]=G_114_0;
   assign c[116]=G_115_0;
   assign c[117]=G_116_0;
   assign c[118]=G_117_0;
   assign c[119]=G_118_0;
   assign c[120]=G_119_0;
   assign c[121]=G_120_0;

   assign c[122]=G_121_0;
   assign c[123]=G_122_0;
   assign c[124]=G_123_0;
   assign c[125]=G_124_0;
   assign c[126]=G_125_0;
   assign c[127]=G_126_0;
   assign c[128]=G_127_0;

endmodule // brent_kung_cs



`timescale 1 ns/10 ps
module tb;


 reg 		[63:0]		xrf;
 reg 		[63:0]		y;
 reg 		[63:0]		zrf;
 reg 						rn;
 reg 						rz;
 reg 						rm;
 reg 						rp;
 reg 		[63:0]		earlyres;
 reg 						earlyressel;
 reg 		[1:0]			bypsel;
 reg 						bypplus1;
 reg 						byppostnorm;
 wire 	[63:0]		w;
 wire 	[63:0]		wbypass;
 wire 		 			invalid;
 wire 					overflow;
 wire 					underflow;
 wire 					inexact;

reg [5:0] i;
integer fp;

localparam period = 20;  
fmac UUT(.xrf(xrf), .y(y), .zrf(zrf), .rn(rn), .rz(rz), .rp(rp), .rm(rm),
		.earlyres(earlyres), .earlyressel(earlyressel), .bypsel(bypsel), .bypplus1(bypplus1), .byppostnorm(byppostnorm), 
		.w(w), .wbypass(wbypass), .invalid(invalid), .overflow(overflow), .underflow(underflow), .inexact(inexact));


initial 
    begin
fp = $fopen("output","w");
    xrf = 64'hc22000007fffffff;
    y = 64'h24700000ffffffef;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfc00000000011fe;
    y = 64'h3fdfffffffffff03;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'ha83100000007fffe;
    y = 64'h41e0000effffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h001ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h400327ca64d70ec7;
    y = 64'h3ca0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h43e207ffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h3fd0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h3fdfffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h3fe0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc870200000010000;
    y = 64'h3fefffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc00aaa4fd557ef13;
    y = 64'hc3b8917384eb32d0;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hc18aca47203438e2;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h4000000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h47efff0008000000;
    y = 64'hb1dcb0523546117f;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43f000ffffff7fff;
    y = 64'h22300000001fffdf;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h402ff000001fffff;
    y = 64'h40759558e27de226;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h40efdeffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h434fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h7ffc000000000000;
    y = 64'h7fe0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb35e061abc769f3a;
    y = 64'hc078000003fffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h403a793cfb1e2471;
    y = 64'hbff0000100007fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3d1ffffbfe000000;
    y = 64'h216898822a24af3f;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfb00000001bffff;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h37f0000000efffff;
    y = 64'hc3d00007fffffeff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hffefff8000080000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fb00200000000ff;
    y = 64'hc0000000011fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41c0000007ffffff;
    y = 64'h49103fffefffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h407effbfffffffff;
    y = 64'h3e00000040001fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1f00013fffffffe;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc3f00004000001ff;
    y = 64'hc3d00bfffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h403b5ab30b28be12;
    y = 64'hbfdfffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hc1cfffffff87ffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hbfe0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h801ffc000007ffff;
    y = 64'hbfeffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hffe0000005fffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hbfffffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hc000000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc3d09308769f3f51;
    y = 64'hc00fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h402ffffdfefffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hc010000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc01fffffffc00fff;
    y = 64'hc01ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc025e14360f49046;
    y = 64'h412fff0000000003;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h43ee59a2f1155c8b;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fe0000000008fff;
    y = 64'h802ffffff7fffff6;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hffefffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h40401007fffffffe;
    y = 64'hfff0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'hc0045abb4860cbf3;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0000000000000000;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbffffffec0000000;
    y = 64'hc000000000003eff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h48000000004001ff;
    y = 64'h41f331de979ac49e;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3d0fffffbff7ffff;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43d3ffffff000000;
    y = 64'h3caffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h7ffc000000000000;
    y = 64'h43dfff8004000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbcaffe0000000008;
    y = 64'h3fd00008000000ff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h404ffbfffffffffc;
    y = 64'hc34ffff8003fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43e0000000000082;
    y = 64'h3db000003ffffeff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1d004000ffffffe;
    y = 64'h4000000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc00fffffc000007e;
    y = 64'hc02ffffdfffffbff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h409dfffbffffffff;
    y = 64'h4010000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc120000003ffffe0;
    y = 64'hc06000fffbffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fd1f7ffffffffff;
    y = 64'hc01000001dffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h2e0fefdfffffffff;
    y = 64'h4030000020000040;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43c0000803ffffff;
    y = 64'h3fcfffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0afffffbffffdfe;
    y = 64'h3fc07ffdffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0fffffffeffffee;
    y = 64'h55139bb9349e058c;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41ffdbaf18ce06bd;
    y = 64'h8010000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0e1000000080000;
    y = 64'h801ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fbffffff0000007;
    y = 64'hc807dfffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc357b53537b96da5;
    y = 64'hbfd0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h401fffffffffffff;
    y = 64'hffebff8000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc7eff77bf2b59c3c;
    y = 64'hbfe0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h380c3f72cc3dec98;
    y = 64'hc3fffffffbffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb8e0000003fbffff;
    y = 64'hc503f4d44f4bf888;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3f3ffffc001fffff;
    y = 64'hc000000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc340002000004000;
    y = 64'hc0db3367e0423019;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h4f60000801ffffff;
    y = 64'h41c07fe000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1ffffffbfefffff;
    y = 64'hc340000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h404fff7fffffff7f;
    y = 64'h48ab7e2aad4ec686;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h7ffc000000000000;
    y = 64'hffefffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41e189ea1a6fff97;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3ff0ee9046c9330f;
    y = 64'h8479e1e79766e02b;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hd2f805130a8c11df;
    y = 64'h43effffdfdfffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h4f1fffbfffe00000;
    y = 64'hbcd02000000007ff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbe70000077ffffff;
    y = 64'hc1efffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41e1ffffbffffffe;
    y = 64'h3caffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3bbd976272fb1d2a;
    y = 64'hc06ffff80007fffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h434fff01ffffffff;
    y = 64'h403dfeffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbe6fff7fffffffff;
    y = 64'h3feffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41d007ff80000000;
    y = 64'h41f0fffffffc0000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hffeef7a206029708;
    y = 64'hbdcfa4109a3a5b22;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3b6ffffffeffffc0;
    y = 64'h3c7ffffe003ffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1d1ffffffbfffff;
    y = 64'hbfcffffefffff800;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h2030000000000090;
    y = 64'hc05e2e90015c47a1;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbbf000000007efff;
    y = 64'h001fe0000007fffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41cae866712069f4;
    y = 64'hc02fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfce1e32ccf56348;
    y = 64'h3ca1f66d4c8eeef3;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hffedfffff0000000;
    y = 64'hffeffff000000800;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h37effffc3ffffffe;
    y = 64'hbca0fffffffffffd;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbc950a021bf9dee1;
    y = 64'h3db0001fffdffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hfd4fffffdfffffef;
    y = 64'h41cffffdffffffef;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfc00000004007ff;
    y = 64'hbcafffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc009130b80fe8274;
    y = 64'hb811571307061a38;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0600000ffffffdf;
    y = 64'h7feda1b8c591f9c6;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1e4af3f8d45e031;
    y = 64'h3ca0020002000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3800008100000000;
    y = 64'hb810000020000080;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h372ff00000003fff;
    y = 64'h7fe000fdfffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h47d00021fffffffe;
    y = 64'hc00fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfbc9ea0c2b4884b;
    y = 64'h43f4a552574073d5;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbf1fe0000000ffff;
    y = 64'hc01ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41ffffffff7ffffb;
    y = 64'h0027ffffffffeffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc7e040000fffffff;
    y = 64'hffe0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h7ffc000000000000;
    y = 64'h3fe0000ffffff7ff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1effc1fffffffff;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0d000000001ffbf;
    y = 64'hc03ba46e644e4e9c;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc4500000005fffff;
    y = 64'hc03a20ab4de47fc9;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h400e00000000007e;
    y = 64'h001fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h45a01fffff7fffff;
    y = 64'hc3c0020200000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3e8ff800000000ff;
    y = 64'h3caffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbe004000000007fe;
    y = 64'h3fdffff7ff7fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb11000007ffffe00;
    y = 64'h3fe0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb80cef50bd17db40;
    y = 64'hc05fffc00000000e;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3d4000ffffffffff;
    y = 64'h3d47f68d8eb6b9a4;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hffe3fffffffffffb;
    y = 64'hc03dc3321aaa5380;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3ca3fffffffffeff;
    y = 64'hbf02ffafb4e9241d;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h53598c812c3c39dd;
    y = 64'h3f20000100fffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc3dffffff8000001;
    y = 64'h3fe0020000003ffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h7ba00800003fffff;
    y = 64'h3ff9a9a129c791b3;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc3d0000fffffffef;
    y = 64'h7fe0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc34f80001fffffff;
    y = 64'hb7fffffe0007ffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000001ff8;
    y = 64'h4800020000010000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h2c4c0000003fffff;
    y = 64'h230ffffc00400000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h381fffffffbff7fe;
    y = 64'h8010000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h802d3018ea8c241d;
    y = 64'hc007fdffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43e047fffffffffe;
    y = 64'h4000003ffdfffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc000005fffffffff;
    y = 64'h403ffffffff00002;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fc8b60e46a80f6d;
    y = 64'hbfdffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbd5fdffdffffffff;
    y = 64'h5644b72ace1bbb6b;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb80010001fffffff;
    y = 64'h40e01ffffff7fffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h407000003ffbfffe;
    y = 64'h38042862fe8e3368;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbf8ffbfff7ffffff;
    y = 64'hc00fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbcafc000003fffff;
    y = 64'hc010000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h47eddf042473ef08;
    y = 64'hb7e00000fe000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3fbfffff7fffffef;
    y = 64'hc340ffffffffffbf;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc02f8000000007ff;
    y = 64'hffe0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h002f37ebf6c8eaec;
    y = 64'hc08be464f4c81c69;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc00e800000000000;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h0000000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbfffc00000000003;
    y = 64'h391001ffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1db54446247aa52;
    y = 64'hbfcc001fffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hc0392c59c8e48f37;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hc0000800000001ff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hc1d0000004000fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h4030040000200000;
    y = 64'h0017055f48beeff5;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbc7000000000ffee;
    y = 64'hc1e0001100000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc040000000007fff;
    y = 64'hc3b2a6c91c557f56;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41ffffffff003fff;
    y = 64'hc3b0000007ffffee;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h21900001dfffffff;
    y = 64'hbf20000017fffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0029954d0f0df5b3;
    y = 64'h41e00000000003ff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb810000020000001;
    y = 64'h47ffdfffffffff80;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hffeffff800007fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h4010000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbf700000000100ff;
    y = 64'h401fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h37feffffffffffff;
    y = 64'h47ef8000000fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb80f800001fffffe;
    y = 64'h44e00000ffff7fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h434ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41ffffdfffff8000;
    y = 64'h7fe0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb80a16ad02c87cd3;
    y = 64'h380fffffffffe7fe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h47f0fffffffffffb;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h41ffffffffbfff7f;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h8000000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc3d00001000001ff;
    y = 64'hb7f60cb3edb38762;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h8010000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43c0007fffdfffff;
    y = 64'h801ffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc7efffffdffffbff;
    y = 64'hbca0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hc11ff00000000003;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hbfd0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc0ffffffffeffffe;
    y = 64'hbfdfffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h6f7000000001fdff;
    y = 64'h1510010000000fff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h37f002000000000f;
    y = 64'hb1effcfffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hcc3050bc013d7cd7;
    y = 64'hbff0000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h87fff0000000fffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hbffffffffffffffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h43effbfffffff7ff;
    y = 64'h7fefffffff801ffe;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc015834380f2b995;
    y = 64'h3f9fff0000000400;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h41dfffffc0001000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'hc01fffffffffffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h41e010000000001f;
    y = 64'hc5b04000000fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h3b40018000000000;
    y = 64'h3ea0400000000100;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h4cdffeffff7fffff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h16dff0001ffffffe;
    y = 64'h3fb500ae0796659d;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hb7e003ffffffff7f;
    y = 64'hdeafffffeffffffd;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h406000001fffbfff;
    y = 64'h3f20020000080000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h0010000000000000;
    y = 64'h7ffc000000000000;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h439fbffffffbffff;
    y = 64'hbf8454fd38ef0ba0;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hc1c000000200007e;
    y = 64'hbf000001ffffffbf;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h480000000008fffe;
    y = 64'h001637e790e69de2;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'hbffffffc000003fe;
    y = 64'h3ca0000000000001;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
    xrf = 64'h6b4848a9a8c0dcd5;
    y = 64'h480ffffffffbdfff;
    zrf = 64'h0000000000000000;
    rn = 1;
    rz = 0;
    rm = 0;
    rp = 0;
    earlyres = 64'b0;
    earlyressel = 0;
    bypsel= 2'b0;
    bypplus1 = 0;
    byppostnorm = 0;
#10
	$fwrite(fp, "%h %h %h\n",xrf,y,w);
	$stop;
	end
endmodule
../../../config/rv64gc/coverage.svh
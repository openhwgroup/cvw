typedef enum logic[3:0] {BP_TWOBIT, BP_GSHARE, BP_GLOBAL, BP_GSHARE_BASIC, 
               BP_GLOBAL_BASIC, BP_LOCAL_BASIC, BP_LOCAL_AHEAD, BP_LOCAL_REPAIR} BranchPredictorType;


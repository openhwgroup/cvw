`define LIB SKY130

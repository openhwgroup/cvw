module sbtm_a2 (input  logic [6:0] a,
		output logic [12:0] y);
   always_comb
     case(a)
       7'b0000000: y = 13'b1111111110001;
       7'b0000001: y = 13'b1111111010001;
       7'b0000010: y = 13'b1111110110010;
       7'b0000011: y = 13'b1111110010011;
       7'b0000100: y = 13'b1111101110101;
       7'b0000101: y = 13'b1111101010110;
       7'b0000110: y = 13'b1111100111001;
       7'b0000111: y = 13'b1111100011011;
       7'b0001000: y = 13'b1111011111110;
       7'b0001001: y = 13'b1111011100001;
       7'b0001010: y = 13'b1111011000100;
       7'b0001011: y = 13'b1111010101000;
       7'b0001100: y = 13'b1111010001100;
       7'b0001101: y = 13'b1111001110000;
       7'b0001110: y = 13'b1111001010101;
       7'b0001111: y = 13'b1111000111010;
       7'b0010000: y = 13'b1111000011111;
       7'b0010001: y = 13'b1111000000100;
       7'b0010010: y = 13'b1110111101010;
       7'b0010011: y = 13'b1110111010000;
       7'b0010100: y = 13'b1110110110110;
       7'b0010101: y = 13'b1110110011101;
       7'b0010110: y = 13'b1110110000100;
       7'b0010111: y = 13'b1110101101011;
       7'b0011000: y = 13'b1110101010010;
       7'b0011001: y = 13'b1110100111001;
       7'b0011010: y = 13'b1110100100001;
       7'b0011011: y = 13'b1110100001001;
       7'b0011100: y = 13'b1110011110001;
       7'b0011101: y = 13'b1110011011010;
       7'b0011110: y = 13'b1110011000010;
       7'b0011111: y = 13'b1110010101011;
       7'b0100000: y = 13'b1110010010100;
       7'b0100001: y = 13'b1110001111110;
       7'b0100010: y = 13'b1110001100111;
       7'b0100011: y = 13'b1110001010001;
       7'b0100100: y = 13'b1110000111011;
       7'b0100101: y = 13'b1110000100101;
       7'b0100110: y = 13'b1110000001111;
       7'b0100111: y = 13'b1101111111010;
       7'b0101000: y = 13'b1101111100101;
       7'b0101001: y = 13'b1101111010000;
       7'b0101010: y = 13'b1101110111011;
       7'b0101011: y = 13'b1101110100110;
       7'b0101100: y = 13'b1101110010001;
       7'b0101101: y = 13'b1101101111101;
       7'b0101110: y = 13'b1101101101001;
       7'b0101111: y = 13'b1101101010101;
       7'b0110000: y = 13'b1101101000001;
       7'b0110001: y = 13'b1101100101101;
       7'b0110010: y = 13'b1101100011010;
       7'b0110011: y = 13'b1101100000110;
       7'b0110100: y = 13'b1101011110011;
       7'b0110101: y = 13'b1101011100000;
       7'b0110110: y = 13'b1101011001101;
       7'b0110111: y = 13'b1101010111010;
       7'b0111000: y = 13'b1101010101000;
       7'b0111001: y = 13'b1101010010101;
       7'b0111010: y = 13'b1101010000011;
       7'b0111011: y = 13'b1101001110001;
       7'b0111100: y = 13'b1101001011111;
       7'b0111101: y = 13'b1101001001101;
       7'b0111110: y = 13'b1101000111100;
       7'b0111111: y = 13'b1101000101010;
       7'b1000000: y = 13'b1101000011001;
       7'b1000001: y = 13'b1101000000111;
       7'b1000010: y = 13'b1100111110110;
       7'b1000011: y = 13'b1100111100101;
       7'b1000100: y = 13'b1100111010100;
       7'b1000101: y = 13'b1100111000011;
       7'b1000110: y = 13'b1100110110011;
       7'b1000111: y = 13'b1100110100010;
       7'b1001000: y = 13'b1100110010010;
       7'b1001001: y = 13'b1100110000010;
       7'b1001010: y = 13'b1100101110010;
       7'b1001011: y = 13'b1100101100001;
       7'b1001100: y = 13'b1100101010010;
       7'b1001101: y = 13'b1100101000010;
       7'b1001110: y = 13'b1100100110010;
       7'b1001111: y = 13'b1100100100011;
       7'b1010000: y = 13'b1100100010011;
       7'b1010001: y = 13'b1100100000100;
       7'b1010010: y = 13'b1100011110101;
       7'b1010011: y = 13'b1100011100101;
       7'b1010100: y = 13'b1100011010110;
       7'b1010101: y = 13'b1100011000111;
       7'b1010110: y = 13'b1100010111001;
       7'b1010111: y = 13'b1100010101010;
       7'b1011000: y = 13'b1100010011011;
       7'b1011001: y = 13'b1100010001101;
       7'b1011010: y = 13'b1100001111110;
       7'b1011011: y = 13'b1100001110000;
       7'b1011100: y = 13'b1100001100010;
       7'b1011101: y = 13'b1100001010100;
       7'b1011110: y = 13'b1100001000110;
       7'b1011111: y = 13'b1100000111000;
       7'b1100000: y = 13'b1100000101010;
       7'b1100001: y = 13'b1100000011100;
       7'b1100010: y = 13'b1100000001111;
       7'b1100011: y = 13'b1100000000001;
       7'b1100100: y = 13'b1011111110100;
       7'b1100101: y = 13'b1011111100110;
       7'b1100110: y = 13'b1011111011001;
       7'b1100111: y = 13'b1011111001100;
       7'b1101000: y = 13'b1011110111111;
       7'b1101001: y = 13'b1011110110010;
       7'b1101010: y = 13'b1011110100101;
       7'b1101011: y = 13'b1011110011000;
       7'b1101100: y = 13'b1011110001011;
       7'b1101101: y = 13'b1011101111110;
       7'b1101110: y = 13'b1011101110010;
       7'b1101111: y = 13'b1011101100101;
       7'b1110000: y = 13'b1011101011001;
       7'b1110001: y = 13'b1011101001100;
       7'b1110010: y = 13'b1011101000000;
       7'b1110011: y = 13'b1011100110100;
       7'b1110100: y = 13'b1011100101000;
       7'b1110101: y = 13'b1011100011100;
       7'b1110110: y = 13'b1011100010000;
       7'b1110111: y = 13'b1011100000100;
       7'b1111000: y = 13'b1011011111000;
       7'b1111001: y = 13'b1011011101100;
       7'b1111010: y = 13'b1011011100000;
       7'b1111011: y = 13'b1011011010101;
       7'b1111100: y = 13'b1011011001001;
       7'b1111101: y = 13'b1011010111101;
       7'b1111110: y = 13'b1011010110010;
       7'b1111111: y = 13'b1011010100111;	    
       default: y = 13'bxxxxxxxxxxxxx;
     endcase // case (a)
    
endmodule // sbtm_a0

    
    
    
///////////////////////////////////////////
// tests.vh
//
// Written: David_Harris@hmc.edu 7 October 2021
// Modified: 
//
// Purpose: List of tests to apply
// 
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define IMPERASTEST   "0"
`define RISCVARCHTEST "1"
`define WALLYTEST "2"
`define MYIMPERASTEST   "3"
`define COREMARK "4"
`define EMBENCH "5"
`define CUSTOM "6"
// *** remove MYIMPERASTEST cases when ported 

string tvpaths[] = '{
    "../addins/imperas-riscv-tests/work/",
    "../tests/riscof/work/riscv-arch-test/",
    "../tests/riscof/work/wally-riscv-arch-test/",
    "../tests/imperas-riscv-tests/work/",
    "../benchmarks/coremark/work/",
    "../addins/embench-iot/",
    "../tests/custom/work/"
    };

  string coremark[] = '{
    `COREMARK,
    "coremark.bare.riscv"
  };

  string embench[] = '{
    `EMBENCH,
    "bd_speedopt_speed/src/nsichneu/nsichneu",
    "bd_speedopt_speed/src/cubic/cubic", // cubic is likely going to removed when embench 2.0 launches
    "bd_speedopt_speed/src/aha-mont64/aha-mont64",
    "bd_speedopt_speed/src/crc32/crc32",
    "bd_speedopt_speed/src/cubic/cubic", // cubic is likely going to removed when embench 2.0 launches
    "bd_speedopt_speed/src/edn/edn",
    "bd_speedopt_speed/src/huffbench/huffbench",
    "bd_speedopt_speed/src/matmult-int/matmult-int",
    // "bd_speedopt_speed/src/md5sum/md5sum", //commenting out tests from embench 2.0. When embench 2.0 launches stabilty, add these tests back
    "bd_speedopt_speed/src/minver/minver",
    "bd_speedopt_speed/src/nettle-aes/nettle-aes",
    "bd_speedopt_speed/src/nettle-sha256/nettle-sha256",
    "bd_speedopt_speed/src/nbody/nbody",
    "bd_speedopt_speed/src/picojpeg/picojpeg",
    // "bd_speedopt_speed/src/primecount/primecount",
    "bd_speedopt_speed/src/qrduino/qrduino",
    "bd_speedopt_speed/src/sglib-combined/sglib-combined",
    "bd_speedopt_speed/src/slre/slre",
    "bd_speedopt_speed/src/st/st",
    "bd_speedopt_speed/src/statemate/statemate",
    // "bd_speedopt_speed/src/tarfind/tarfind",
    "bd_speedopt_speed/src/ud/ud",
    "bd_speedopt_speed/src/wikisort/wikisort",
    "bd_sizeopt_speed/src/aha-mont64/aha-mont64",
    "bd_sizeopt_speed/src/crc32/crc32",
    "bd_sizeopt_speed/src/cubic/cubic",
    "bd_sizeopt_speed/src/edn/edn",
    "bd_sizeopt_speed/src/huffbench/huffbench",
    "bd_sizeopt_speed/src/matmult-int/matmult-int",
    // "bd_sizeopt_speed/src/md5sum/md5sum",
    "bd_sizeopt_speed/src/minver/minver",
    "bd_sizeopt_speed/src/nbody/nbody",
    "bd_sizeopt_speed/src/nettle-aes/nettle-aes",
    "bd_sizeopt_speed/src/nettle-sha256/nettle-sha256",
    "bd_sizeopt_speed/src/nsichneu/nsichneu",
    "bd_sizeopt_speed/src/picojpeg/picojpeg",
    // "bd_sizeopt_speed/src/primecount/primecount",
    "bd_sizeopt_speed/src/qrduino/qrduino",
    "bd_sizeopt_speed/src/sglib-combined/sglib-combined",
    "bd_sizeopt_speed/src/slre/slre",
    "bd_sizeopt_speed/src/st/st",
    "bd_sizeopt_speed/src/statemate/statemate",
    // "bd_sizeopt_speed/src/tarfind/tarfind",
    "bd_sizeopt_speed/src/ud/ud",
    "bd_sizeopt_speed/src/wikisort/wikisort"
  };
  
string imperas32f[] = '{
    `IMPERASTEST,
    "rv32i_m/F/FSQRT-S-DYN-RDN-01.S",
    "rv32i_m/F/FADD-S-DYN-RDN-01.S",
    "rv32i_m/F/FADD-S-DYN-RMM-01.S",
    "rv32i_m/F/FADD-S-DYN-RNE-01.S",
    "rv32i_m/F/FADD-S-DYN-RTZ-01.S",
    "rv32i_m/F/FADD-S-DYN-RUP-01.S",
    "rv32i_m/F/FADD-S-RDN-01.S",
    "rv32i_m/F/FADD-S-RMM-01.S",
    "rv32i_m/F/FADD-S-RNE-01.S",
    "rv32i_m/F/FADD-S-RTZ-01.S",
    "rv32i_m/F/FADD-S-RUP-01.S",
    "rv32i_m/F/FCLASS-S-01.S",
    "rv32i_m/F/FCVT-S-W-DYN-RDN-01.S",
    "rv32i_m/F/FCVT-S-W-DYN-RMM-01.S",
    "rv32i_m/F/FCVT-S-W-DYN-RNE-01.S",
    "rv32i_m/F/FCVT-S-W-DYN-RTZ-01.S",
    "rv32i_m/F/FCVT-S-W-DYN-RUP-01.S",
    "rv32i_m/F/FCVT-S-W-RDN-01.S",
    "rv32i_m/F/FCVT-S-W-RMM-01.S",
    "rv32i_m/F/FCVT-S-W-RNE-01.S",
    "rv32i_m/F/FCVT-S-W-RTZ-01.S",
    "rv32i_m/F/FCVT-S-W-RUP-01.S",
    "rv32i_m/F/FCVT-S-WU-DYN-RDN-01.S",
    "rv32i_m/F/FCVT-S-WU-DYN-RMM-01.S",
    "rv32i_m/F/FCVT-S-WU-DYN-RNE-01.S",
    "rv32i_m/F/FCVT-S-WU-DYN-RTZ-01.S",
    "rv32i_m/F/FCVT-S-WU-DYN-RUP-01.S",
    "rv32i_m/F/FCVT-S-WU-RDN-01.S",
    "rv32i_m/F/FCVT-S-WU-RMM-01.S",
    "rv32i_m/F/FCVT-S-WU-RNE-01.S",
    "rv32i_m/F/FCVT-S-WU-RTZ-01.S",
    "rv32i_m/F/FCVT-S-WU-RUP-01.S",
    "rv32i_m/F/FCVT-W-S-DYN-RDN-01.S",
    "rv32i_m/F/FCVT-W-S-DYN-RMM-01.S",
    "rv32i_m/F/FCVT-W-S-DYN-RNE-01.S",
    "rv32i_m/F/FCVT-W-S-DYN-RTZ-01.S",
    "rv32i_m/F/FCVT-W-S-DYN-RUP-01.S",
    "rv32i_m/F/FCVT-W-S-RDN-01.S",
    "rv32i_m/F/FCVT-W-S-RMM-01.S",
    "rv32i_m/F/FCVT-W-S-RNE-01.S",
    "rv32i_m/F/FCVT-W-S-RTZ-01.S",
    "rv32i_m/F/FCVT-W-S-RUP-01.S",
    "rv32i_m/F/FCVT-WU-S-DYN-RDN-01.S",
    "rv32i_m/F/FCVT-WU-S-DYN-RMM-01.S",
    "rv32i_m/F/FCVT-WU-S-DYN-RNE-01.S",
    "rv32i_m/F/FCVT-WU-S-DYN-RTZ-01.S",
    "rv32i_m/F/FCVT-WU-S-DYN-RUP-01.S",
    "rv32i_m/F/FCVT-WU-S-RDN-01.S",
    "rv32i_m/F/FCVT-WU-S-RMM-01.S",
    "rv32i_m/F/FCVT-WU-S-RNE-01.S",
    "rv32i_m/F/FCVT-WU-S-RTZ-01.S",
    "rv32i_m/F/FCVT-WU-S-RUP-01.S",
    "rv32i_m/F/FDIV-S-DYN-RDN-01.S",
    "rv32i_m/F/FDIV-S-DYN-RMM-01.S",
    "rv32i_m/F/FDIV-S-DYN-RNE-01.S",
    "rv32i_m/F/FDIV-S-DYN-RTZ-01.S",
    "rv32i_m/F/FDIV-S-DYN-RUP-01.S",
    "rv32i_m/F/FDIV-S-RDN-01.S",
    "rv32i_m/F/FDIV-S-RMM-01.S",
    "rv32i_m/F/FDIV-S-RNE-01.S",
    "rv32i_m/F/FDIV-S-RTZ-01.S",
    "rv32i_m/F/FDIV-S-RUP-01.S",
    "rv32i_m/F/FEQ-S-01.S",
    "rv32i_m/F/FLE-S-01.S",
    "rv32i_m/F/FLT-S-01.S",
    "rv32i_m/F/FLW-01.S",
    "rv32i_m/F/FMADD-S-DYN-RDN-01.S",
    "rv32i_m/F/FMADD-S-DYN-RMM-01.S",
    "rv32i_m/F/FMADD-S-DYN-RNE-01.S",
    "rv32i_m/F/FMADD-S-DYN-RTZ-01.S",
    "rv32i_m/F/FMADD-S-DYN-RUP-01.S",
    "rv32i_m/F/FMADD-S-RDN-01.S",
    "rv32i_m/F/FMADD-S-RMM-01.S",
    "rv32i_m/F/FMADD-S-RNE-01.S",
    "rv32i_m/F/FMADD-S-RTZ-01.S",
    "rv32i_m/F/FMADD-S-RUP-01.S",
    "rv32i_m/F/FMAX-S-01.S",
    "rv32i_m/F/FMIN-S-01.S",
    "rv32i_m/F/FMSUB-S-DYN-RDN-01.S",
    "rv32i_m/F/FMSUB-S-DYN-RMM-01.S",
    "rv32i_m/F/FMSUB-S-DYN-RNE-01.S",
    "rv32i_m/F/FMSUB-S-DYN-RTZ-01.S",
    "rv32i_m/F/FMSUB-S-DYN-RUP-01.S",
    "rv32i_m/F/FMSUB-S-RDN-01.S",
    "rv32i_m/F/FMSUB-S-RMM-01.S",
    "rv32i_m/F/FMSUB-S-RNE-01.S",
    "rv32i_m/F/FMSUB-S-RTZ-01.S",
    "rv32i_m/F/FMSUB-S-RUP-01.S",
    "rv32i_m/F/FMUL-S-DYN-RDN-01.S",
    "rv32i_m/F/FMUL-S-DYN-RMM-01.S",
    "rv32i_m/F/FMUL-S-DYN-RNE-01.S",
    "rv32i_m/F/FMUL-S-DYN-RTZ-01.S",
    "rv32i_m/F/FMUL-S-DYN-RUP-01.S",
    "rv32i_m/F/FMUL-S-RDN-01.S",
    "rv32i_m/F/FMUL-S-RMM-01.S",
    "rv32i_m/F/FMUL-S-RNE-01.S",
    "rv32i_m/F/FMUL-S-RTZ-01.S",
    "rv32i_m/F/FMUL-S-RUP-01.S",
    "rv32i_m/F/FMV-W-X-01.S",
    "rv32i_m/F/FMV-X-W-01.S",
    "rv32i_m/F/FNMADD-S-DYN-RDN-01.S",
    "rv32i_m/F/FNMADD-S-DYN-RMM-01.S",
    "rv32i_m/F/FNMADD-S-DYN-RNE-01.S",
    "rv32i_m/F/FNMADD-S-DYN-RTZ-01.S",
    "rv32i_m/F/FNMADD-S-DYN-RUP-01.S",
    "rv32i_m/F/FNMADD-S-RDN-01.S",
    "rv32i_m/F/FNMADD-S-RMM-01.S",
    "rv32i_m/F/FNMADD-S-RNE-01.S",
    "rv32i_m/F/FNMADD-S-RTZ-01.S",
    "rv32i_m/F/FNMADD-S-RUP-01.S",
    "rv32i_m/F/FNMSUB-S-DYN-RDN-01.S",
    "rv32i_m/F/FNMSUB-S-DYN-RMM-01.S",
    "rv32i_m/F/FNMSUB-S-DYN-RNE-01.S",
    "rv32i_m/F/FNMSUB-S-DYN-RTZ-01.S",
    "rv32i_m/F/FNMSUB-S-DYN-RUP-01.S",
    "rv32i_m/F/FNMSUB-S-RDN-01.S",
    "rv32i_m/F/FNMSUB-S-RMM-01.S",
    "rv32i_m/F/FNMSUB-S-RNE-01.S",
    "rv32i_m/F/FNMSUB-S-RTZ-01.S",
    "rv32i_m/F/FNMSUB-S-RUP-01.S",
    "rv32i_m/F/FSGNJN-S-01.S",
    "rv32i_m/F/FSGNJ-S-01.S",
    "rv32i_m/F/FSGNJX-S-01.S",
    "rv32i_m/F/FSQRT-S-DYN-RDN-01.S",
    "rv32i_m/F/FSQRT-S-DYN-RMM-01.S",
    "rv32i_m/F/FSQRT-S-DYN-RNE-01.S",
    "rv32i_m/F/FSQRT-S-DYN-RTZ-01.S",
    "rv32i_m/F/FSQRT-S-DYN-RUP-01.S",
    "rv32i_m/F/FSQRT-S-RDN-01.S",
    "rv32i_m/F/FSQRT-S-RMM-01.S",
    "rv32i_m/F/FSQRT-S-RNE-01.S",
    "rv32i_m/F/FSQRT-S-RTZ-01.S",
    "rv32i_m/F/FSQRT-S-RUP-01.S",
    "rv32i_m/F/FSUB-S-DYN-RDN-01.S",
    "rv32i_m/F/FSUB-S-DYN-RMM-01.S",
    "rv32i_m/F/FSUB-S-DYN-RNE-01.S",
    "rv32i_m/F/FSUB-S-DYN-RTZ-01.S",
    "rv32i_m/F/FSUB-S-DYN-RUP-01.S",
    "rv32i_m/F/FSUB-S-RDN-01.S",
    "rv32i_m/F/FSUB-S-RMM-01.S",
    "rv32i_m/F/FSUB-S-RNE-01.S",
    "rv32i_m/F/FSUB-S-RTZ-01.S",
    "rv32i_m/F/FSUB-S-RUP-01.S",
    "rv32i_m/F/FSW-01.S"
  };

  string imperas64f[] = '{
    `IMPERASTEST,
    "rv64i_m/F/FADD-S-DYN-RDN-01.S",
    "rv64i_m/F/FADD-S-DYN-RMM-01.S",
    "rv64i_m/F/FADD-S-DYN-RNE-01.S",
    "rv64i_m/F/FADD-S-DYN-RTZ-01.S",
    "rv64i_m/F/FADD-S-DYN-RUP-01.S",
    "rv64i_m/F/FADD-S-RDN-01.S",
    "rv64i_m/F/FADD-S-RMM-01.S",
    "rv64i_m/F/FADD-S-RNE-01.S",
    "rv64i_m/F/FADD-S-RTZ-01.S",
    "rv64i_m/F/FADD-S-RUP-01.S",
    "rv64i_m/F/FCLASS-S-01.S",
    "rv64i_m/F/FCVT-L-S-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-L-S-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-L-S-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-L-S-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-L-S-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-L-S-RDN-01.S",
    "rv64i_m/F/FCVT-L-S-RMM-01.S",
    "rv64i_m/F/FCVT-L-S-RNE-01.S",
    "rv64i_m/F/FCVT-L-S-RTZ-01.S",
    "rv64i_m/F/FCVT-L-S-RUP-01.S",
    "rv64i_m/F/FCVT-LU-S-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-LU-S-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-LU-S-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-LU-S-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-LU-S-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-LU-S-RDN-01.S",
    "rv64i_m/F/FCVT-LU-S-RMM-01.S",
    "rv64i_m/F/FCVT-LU-S-RNE-01.S",
    "rv64i_m/F/FCVT-LU-S-RTZ-01.S",
    "rv64i_m/F/FCVT-LU-S-RUP-01.S",
    "rv64i_m/F/FCVT-S-L-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-S-L-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-S-L-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-S-L-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-S-L-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-S-L-RDN-01.S",
    "rv64i_m/F/FCVT-S-L-RMM-01.S",
    "rv64i_m/F/FCVT-S-L-RNE-01.S",
    "rv64i_m/F/FCVT-S-L-RTZ-01.S",
    "rv64i_m/F/FCVT-S-L-RUP-01.S",
    "rv64i_m/F/FCVT-S-LU-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-S-LU-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-S-LU-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-S-LU-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-S-LU-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-S-LU-RDN-01.S",
    "rv64i_m/F/FCVT-S-LU-RMM-01.S",
    "rv64i_m/F/FCVT-S-LU-RNE-01.S",
    "rv64i_m/F/FCVT-S-LU-RTZ-01.S",
    "rv64i_m/F/FCVT-S-LU-RUP-01.S",
    "rv64i_m/F/FCVT-S-W-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-S-W-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-S-W-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-S-W-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-S-W-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-S-W-RDN-01.S",
    "rv64i_m/F/FCVT-S-W-RMM-01.S",
    "rv64i_m/F/FCVT-S-W-RNE-01.S",
    "rv64i_m/F/FCVT-S-W-RTZ-01.S",
    "rv64i_m/F/FCVT-S-W-RUP-01.S",
    "rv64i_m/F/FCVT-S-WU-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-S-WU-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-S-WU-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-S-WU-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-S-WU-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-S-WU-RDN-01.S",
    "rv64i_m/F/FCVT-S-WU-RMM-01.S",
    "rv64i_m/F/FCVT-S-WU-RNE-01.S",
    "rv64i_m/F/FCVT-S-WU-RTZ-01.S",
    "rv64i_m/F/FCVT-S-WU-RUP-01.S",
    "rv64i_m/F/FCVT-W-S-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-W-S-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-W-S-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-W-S-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-W-S-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-W-S-RDN-01.S",
    "rv64i_m/F/FCVT-W-S-RMM-01.S",
    "rv64i_m/F/FCVT-W-S-RNE-01.S",
    "rv64i_m/F/FCVT-W-S-RTZ-01.S",
    "rv64i_m/F/FCVT-W-S-RUP-01.S",
    "rv64i_m/F/FCVT-WU-S-DYN-RDN-01.S",
    "rv64i_m/F/FCVT-WU-S-DYN-RMM-01.S",
    "rv64i_m/F/FCVT-WU-S-DYN-RNE-01.S",
    "rv64i_m/F/FCVT-WU-S-DYN-RTZ-01.S",
    "rv64i_m/F/FCVT-WU-S-DYN-RUP-01.S",
    "rv64i_m/F/FCVT-WU-S-RDN-01.S",
    "rv64i_m/F/FCVT-WU-S-RMM-01.S",
    "rv64i_m/F/FCVT-WU-S-RNE-01.S",
    "rv64i_m/F/FCVT-WU-S-RTZ-01.S",
    "rv64i_m/F/FCVT-WU-S-RUP-01.S",
    "rv64i_m/F/FDIV-S-DYN-RDN-01.S",
    "rv64i_m/F/FDIV-S-DYN-RMM-01.S",
    "rv64i_m/F/FDIV-S-DYN-RNE-01.S",
    "rv64i_m/F/FDIV-S-DYN-RTZ-01.S",
    "rv64i_m/F/FDIV-S-DYN-RUP-01.S",
    "rv64i_m/F/FDIV-S-RDN-01.S",
    "rv64i_m/F/FDIV-S-RMM-01.S",
    "rv64i_m/F/FDIV-S-RNE-01.S",
    "rv64i_m/F/FDIV-S-RTZ-01.S",
    "rv64i_m/F/FDIV-S-RUP-01.S",
    "rv64i_m/F/FEQ-S-01.S",
    "rv64i_m/F/FLE-S-01.S",
    "rv64i_m/F/FLT-S-01.S",
    "rv64i_m/F/FLW-01.S",
    "rv64i_m/F/FMADD-S-DYN-RDN-01.S",
    "rv64i_m/F/FMADD-S-DYN-RMM-01.S",
    "rv64i_m/F/FMADD-S-DYN-RNE-01.S",
    "rv64i_m/F/FMADD-S-DYN-RTZ-01.S",
    "rv64i_m/F/FMADD-S-DYN-RUP-01.S",
    "rv64i_m/F/FMADD-S-RDN-01.S",
    "rv64i_m/F/FMADD-S-RMM-01.S",
    "rv64i_m/F/FMADD-S-RNE-01.S",
    "rv64i_m/F/FMADD-S-RTZ-01.S",
    "rv64i_m/F/FMADD-S-RUP-01.S",
    "rv64i_m/F/FMAX-S-01.S",
    "rv64i_m/F/FMIN-S-01.S",
    "rv64i_m/F/FMSUB-S-DYN-RDN-01.S",
    "rv64i_m/F/FMSUB-S-DYN-RMM-01.S",
    "rv64i_m/F/FMSUB-S-DYN-RNE-01.S",
    "rv64i_m/F/FMSUB-S-DYN-RTZ-01.S",
    "rv64i_m/F/FMSUB-S-DYN-RUP-01.S",
    "rv64i_m/F/FMSUB-S-RDN-01.S",
    "rv64i_m/F/FMSUB-S-RMM-01.S",
    "rv64i_m/F/FMSUB-S-RNE-01.S",
    "rv64i_m/F/FMSUB-S-RTZ-01.S",
    "rv64i_m/F/FMSUB-S-RUP-01.S",
    "rv64i_m/F/FMUL-S-DYN-RDN-01.S",
    "rv64i_m/F/FMUL-S-DYN-RMM-01.S",
    "rv64i_m/F/FMUL-S-DYN-RNE-01.S",
    "rv64i_m/F/FMUL-S-DYN-RTZ-01.S",
    "rv64i_m/F/FMUL-S-DYN-RUP-01.S",
    "rv64i_m/F/FMUL-S-RDN-01.S",
    "rv64i_m/F/FMUL-S-RMM-01.S",
    "rv64i_m/F/FMUL-S-RNE-01.S",
    "rv64i_m/F/FMUL-S-RTZ-01.S",
    "rv64i_m/F/FMUL-S-RUP-01.S",
    "rv64i_m/F/FMV-W-X-01.S",
    "rv64i_m/F/FMV-X-W-01.S",
    "rv64i_m/F/FNMADD-S-DYN-RDN-01.S",
    "rv64i_m/F/FNMADD-S-DYN-RMM-01.S",
    "rv64i_m/F/FNMADD-S-DYN-RNE-01.S",
    "rv64i_m/F/FNMADD-S-DYN-RTZ-01.S",
    "rv64i_m/F/FNMADD-S-DYN-RUP-01.S",
    "rv64i_m/F/FNMADD-S-RDN-01.S",
    "rv64i_m/F/FNMADD-S-RMM-01.S",
    "rv64i_m/F/FNMADD-S-RNE-01.S",
    "rv64i_m/F/FNMADD-S-RTZ-01.S",
    "rv64i_m/F/FNMADD-S-RUP-01.S",
    "rv64i_m/F/FNMSUB-S-DYN-RDN-01.S",
    "rv64i_m/F/FNMSUB-S-DYN-RMM-01.S",
    "rv64i_m/F/FNMSUB-S-DYN-RNE-01.S",
    "rv64i_m/F/FNMSUB-S-DYN-RTZ-01.S",
    "rv64i_m/F/FNMSUB-S-DYN-RUP-01.S",
    "rv64i_m/F/FNMSUB-S-RDN-01.S",
    "rv64i_m/F/FNMSUB-S-RMM-01.S",
    "rv64i_m/F/FNMSUB-S-RNE-01.S",
    "rv64i_m/F/FNMSUB-S-RTZ-01.S",
    "rv64i_m/F/FNMSUB-S-RUP-01.S",
    "rv64i_m/F/FSGNJN-S-01.S",
    "rv64i_m/F/FSGNJ-S-01.S",
    "rv64i_m/F/FSGNJX-S-01.S",
    "rv64i_m/F/FSQRT-S-DYN-RDN-01.S",
    "rv64i_m/F/FSQRT-S-DYN-RMM-01.S",
    "rv64i_m/F/FSQRT-S-DYN-RNE-01.S",
    "rv64i_m/F/FSQRT-S-DYN-RTZ-01.S",
    "rv64i_m/F/FSQRT-S-DYN-RUP-01.S",
    "rv64i_m/F/FSQRT-S-RDN-01.S",
    "rv64i_m/F/FSQRT-S-RMM-01.S",
    "rv64i_m/F/FSQRT-S-RNE-01.S",
    "rv64i_m/F/FSQRT-S-RTZ-01.S",
    "rv64i_m/F/FSQRT-S-RUP-01.S",
    "rv64i_m/F/FSUB-S-DYN-RDN-01.S",
    "rv64i_m/F/FSUB-S-DYN-RMM-01.S",
    "rv64i_m/F/FSUB-S-DYN-RNE-01.S",
    "rv64i_m/F/FSUB-S-DYN-RTZ-01.S",
    "rv64i_m/F/FSUB-S-DYN-RUP-01.S",
    "rv64i_m/F/FSUB-S-RDN-01.S",
    "rv64i_m/F/FSUB-S-RMM-01.S",
    "rv64i_m/F/FSUB-S-RNE-01.S",
    "rv64i_m/F/FSUB-S-RTZ-01.S",
    "rv64i_m/F/FSUB-S-RUP-01.S",
    "rv64i_m/F/FSW-01.S"
  };

  string imperas64d[] = '{
    `IMPERASTEST,
    "rv64i_m/D/FADD-D-DYN-RDN-01.S",
    "rv64i_m/D/FADD-D-DYN-RMM-01.S",
    "rv64i_m/D/FADD-D-DYN-RNE-01.S",
    "rv64i_m/D/FADD-D-DYN-RTZ-01.S",
    "rv64i_m/D/FADD-D-DYN-RUP-01.S",
    "rv64i_m/D/FADD-D-RDN-01.S",
    "rv64i_m/D/FADD-D-RMM-01.S",
    "rv64i_m/D/FADD-D-RNE-01.S",
    "rv64i_m/D/FADD-D-RTZ-01.S",
    "rv64i_m/D/FADD-D-RUP-01.S",
    "rv64i_m/D/FCLASS-D-01.S",
    "rv64i_m/D/FCVT-D-L-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-D-L-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-D-L-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-D-L-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-D-L-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-D-L-RDN-01.S",
    "rv64i_m/D/FCVT-D-L-RMM-01.S",
    "rv64i_m/D/FCVT-D-L-RNE-01.S",
    "rv64i_m/D/FCVT-D-L-RTZ-01.S",
    "rv64i_m/D/FCVT-D-L-RUP-01.S",
    "rv64i_m/D/FCVT-D-LU-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-D-LU-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-D-LU-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-D-LU-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-D-LU-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-D-LU-RDN-01.S",
    "rv64i_m/D/FCVT-D-LU-RMM-01.S",
    "rv64i_m/D/FCVT-D-LU-RNE-01.S",
    "rv64i_m/D/FCVT-D-LU-RTZ-01.S",
    "rv64i_m/D/FCVT-D-LU-RUP-01.S",
    "rv64i_m/D/FCVT-D-S-01.S",
    "rv64i_m/D/FCVT-D-W-01.S",
    "rv64i_m/D/FCVT-D-WU-01.S",
    "rv64i_m/D/FCVT-L-D-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-L-D-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-L-D-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-L-D-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-L-D-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-L-D-RDN-01.S",
    "rv64i_m/D/FCVT-L-D-RMM-01.S",
    "rv64i_m/D/FCVT-L-D-RNE-01.S",
    "rv64i_m/D/FCVT-L-D-RTZ-01.S",
    "rv64i_m/D/FCVT-L-D-RUP-01.S",
    "rv64i_m/D/FCVT-LU-D-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-LU-D-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-LU-D-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-LU-D-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-LU-D-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-LU-D-RDN-01.S",
    "rv64i_m/D/FCVT-LU-D-RMM-01.S",
    "rv64i_m/D/FCVT-LU-D-RNE-01.S",
    "rv64i_m/D/FCVT-LU-D-RTZ-01.S",
    "rv64i_m/D/FCVT-LU-D-RUP-01.S",
    "rv64i_m/D/FCVT-S-D-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-S-D-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-S-D-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-S-D-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-S-D-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-S-D-RDN-01.S",
    "rv64i_m/D/FCVT-S-D-RMM-01.S",
    "rv64i_m/D/FCVT-S-D-RNE-01.S",
    "rv64i_m/D/FCVT-S-D-RTZ-01.S",
    "rv64i_m/D/FCVT-S-D-RUP-01.S",
    "rv64i_m/D/FCVT-W-D-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-W-D-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-W-D-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-W-D-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-W-D-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-W-D-RDN-01.S",
    "rv64i_m/D/FCVT-W-D-RMM-01.S",
    "rv64i_m/D/FCVT-W-D-RNE-01.S",
    "rv64i_m/D/FCVT-W-D-RTZ-01.S",
    "rv64i_m/D/FCVT-W-D-RUP-01.S",
    "rv64i_m/D/FCVT-WU-D-DYN-RDN-01.S",
    "rv64i_m/D/FCVT-WU-D-DYN-RMM-01.S",
    "rv64i_m/D/FCVT-WU-D-DYN-RNE-01.S",
    "rv64i_m/D/FCVT-WU-D-DYN-RTZ-01.S",
    "rv64i_m/D/FCVT-WU-D-DYN-RUP-01.S",
    "rv64i_m/D/FCVT-WU-D-RDN-01.S",
    "rv64i_m/D/FCVT-WU-D-RMM-01.S",
    "rv64i_m/D/FCVT-WU-D-RNE-01.S",
    "rv64i_m/D/FCVT-WU-D-RTZ-01.S",
    "rv64i_m/D/FCVT-WU-D-RUP-01.S",
    "rv64i_m/D/FDIV-D-DYN-RDN-01.S",
    "rv64i_m/D/FDIV-D-DYN-RMM-01.S",
    "rv64i_m/D/FDIV-D-DYN-RNE-01.S",
    "rv64i_m/D/FDIV-D-DYN-RTZ-01.S",
    "rv64i_m/D/FDIV-D-DYN-RUP-01.S",
    "rv64i_m/D/FDIV-D-RDN-01.S",
    "rv64i_m/D/FDIV-D-RMM-01.S",
    "rv64i_m/D/FDIV-D-RNE-01.S",
    "rv64i_m/D/FDIV-D-RTZ-01.S",
    "rv64i_m/D/FDIV-D-RUP-01.S",
    "rv64i_m/D/FEQ-D-01.S",
    "rv64i_m/D/FLD-01.S",
    "rv64i_m/D/FLE-D-01.S",
    "rv64i_m/D/FLT-D-01.S",
    "rv64i_m/D/FMADD-D-DYN-RDN-01.S",
    "rv64i_m/D/FMADD-D-DYN-RMM-01.S",
    "rv64i_m/D/FMADD-D-DYN-RNE-01.S",
    "rv64i_m/D/FMADD-D-DYN-RTZ-01.S",
    "rv64i_m/D/FMADD-D-DYN-RUP-01.S",
    "rv64i_m/D/FMADD-D-RDN-01.S",
    "rv64i_m/D/FMADD-D-RMM-01.S",
    "rv64i_m/D/FMADD-D-RNE-01.S",
    "rv64i_m/D/FMADD-D-RTZ-01.S",
    "rv64i_m/D/FMADD-D-RUP-01.S",
    "rv64i_m/D/FMAX-D-01.S",
    "rv64i_m/D/FMIN-D-01.S",
    "rv64i_m/D/FMSUB-D-DYN-RDN-01.S",
    "rv64i_m/D/FMSUB-D-DYN-RMM-01.S",
    "rv64i_m/D/FMSUB-D-DYN-RNE-01.S",
    "rv64i_m/D/FMSUB-D-DYN-RTZ-01.S",
    "rv64i_m/D/FMSUB-D-DYN-RUP-01.S",
    "rv64i_m/D/FMSUB-D-RDN-01.S",
    "rv64i_m/D/FMSUB-D-RMM-01.S",
    "rv64i_m/D/FMSUB-D-RNE-01.S",
    "rv64i_m/D/FMSUB-D-RTZ-01.S",
    "rv64i_m/D/FMSUB-D-RUP-01.S",
    "rv64i_m/D/FMUL-D-DYN-RDN-01.S",
    "rv64i_m/D/FMUL-D-DYN-RMM-01.S",
    "rv64i_m/D/FMUL-D-DYN-RNE-01.S",
    "rv64i_m/D/FMUL-D-DYN-RTZ-01.S",
    "rv64i_m/D/FMUL-D-DYN-RUP-01.S",
    "rv64i_m/D/FMUL-D-RDN-01.S",
    "rv64i_m/D/FMUL-D-RMM-01.S",
    "rv64i_m/D/FMUL-D-RNE-01.S",
    "rv64i_m/D/FMUL-D-RTZ-01.S",
    "rv64i_m/D/FMUL-D-RUP-01.S",
    "rv64i_m/D/FMV-D-X-01.S",
    "rv64i_m/D/FMV-X-D-01.S",
    "rv64i_m/D/FNMADD-D-DYN-RDN-01.S",
    "rv64i_m/D/FNMADD-D-DYN-RMM-01.S",
    "rv64i_m/D/FNMADD-D-DYN-RNE-01.S",
    "rv64i_m/D/FNMADD-D-DYN-RTZ-01.S",
    "rv64i_m/D/FNMADD-D-DYN-RUP-01.S",
    "rv64i_m/D/FNMADD-D-RDN-01.S",
    "rv64i_m/D/FNMADD-D-RMM-01.S",
    "rv64i_m/D/FNMADD-D-RNE-01.S",
    "rv64i_m/D/FNMADD-D-RTZ-01.S",
    "rv64i_m/D/FNMADD-D-RUP-01.S",
    "rv64i_m/D/FNMSUB-D-DYN-RDN-01.S",
    "rv64i_m/D/FNMSUB-D-DYN-RMM-01.S",
    "rv64i_m/D/FNMSUB-D-DYN-RNE-01.S",
    "rv64i_m/D/FNMSUB-D-DYN-RTZ-01.S",
    "rv64i_m/D/FNMSUB-D-DYN-RUP-01.S",
    "rv64i_m/D/FNMSUB-D-RDN-01.S",
    "rv64i_m/D/FNMSUB-D-RMM-01.S",
    "rv64i_m/D/FNMSUB-D-RNE-01.S",
    "rv64i_m/D/FNMSUB-D-RTZ-01.S",
    "rv64i_m/D/FNMSUB-D-RUP-01.S",
    "rv64i_m/D/FSD-01.S",
    "rv64i_m/D/FSGNJ-D-01.S",
    "rv64i_m/D/FSGNJN-D-01.S",
    "rv64i_m/D/FSGNJX-D-01.S",
    "rv64i_m/D/FSQRT-D-DYN-RDN-01.S",
    "rv64i_m/D/FSQRT-D-DYN-RMM-01.S",
    "rv64i_m/D/FSQRT-D-DYN-RNE-01.S",
    "rv64i_m/D/FSQRT-D-DYN-RTZ-01.S",
    "rv64i_m/D/FSQRT-D-DYN-RUP-01.S",
    "rv64i_m/D/FSQRT-D-RDN-01.S",
    "rv64i_m/D/FSQRT-D-RMM-01.S",
    "rv64i_m/D/FSQRT-D-RNE-01.S",
    "rv64i_m/D/FSQRT-D-RTZ-01.S",
    "rv64i_m/D/FSQRT-D-RUP-01.S",
    "rv64i_m/D/FSUB-D-DYN-RDN-01.S",
    "rv64i_m/D/FSUB-D-DYN-RMM-01.S",
    "rv64i_m/D/FSUB-D-DYN-RNE-01.S",
    "rv64i_m/D/FSUB-D-DYN-RTZ-01.S",
    "rv64i_m/D/FSUB-D-DYN-RUP-01.S",
    "rv64i_m/D/FSUB-D-RDN-01.S",
    "rv64i_m/D/FSUB-D-RMM-01.S",
    "rv64i_m/D/FSUB-D-RNE-01.S",
    "rv64i_m/D/FSUB-D-RTZ-01.S",
    "rv64i_m/D/FSUB-D-RUP-01.S"
};

  string imperas64m[] = '{
    `IMPERASTEST,
    "rv64i_m/M/DIV-01.S",
    "rv64i_m/M/DIVU-01.S",
    "rv64i_m/M/DIVUW-01.S",
    "rv64i_m/M/DIVW-01.S",
    "rv64i_m/M/MUL-01.S",
    "rv64i_m/M/MULH-01.S",
    "rv64i_m/M/MULHSU-01.S",
    "rv64i_m/M/MULHU-01.S",
    "rv64i_m/M/MULW-01.S",
    "rv64i_m/M/REM-01.S",
    "rv64i_m/M/REMU-01.S",
    "rv64i_m/M/REMUW-01.S",
    "rv64i_m/M/REMW-01.S"
  };

  string imperas64c[] = '{
    `IMPERASTEST,
    "rv64i_m/C/C-ADD-01.S",
    "rv64i_m/C/C-ADDI-01.S",
    "rv64i_m/C/C-ADDI16SP-01.S",
    "rv64i_m/C/C-ADDI4SPN-01.S",
    "rv64i_m/C/C-ADDIW-01.S",
    "rv64i_m/C/C-ADDW-01.S",
    "rv64i_m/C/C-AND-01.S",
    "rv64i_m/C/C-ANDI-01.S",
    "rv64i_m/C/C-BEQZ-01.S",
    "rv64i_m/C/C-BNEZ-01.S",
    "rv64i_m/C/C-J-01.S",
    "rv64i_m/C/C-JALR-01.S",
    "rv64i_m/C/C-JR-01.S",
    "rv64i_m/C/C-LD-01.S",
    "rv64i_m/C/C-LDSP-01.S",
    "rv64i_m/C/C-LI-01.S",
    "rv64i_m/C/C-LUI-01.S",
    "rv64i_m/C/C-LW-01.S",
    "rv64i_m/C/C-LWSP-01.S",
    "rv64i_m/C/C-MV-01.S",
    "rv64i_m/C/C-OR-01.S",
    "rv64i_m/C/C-SD-01.S",
    "rv64i_m/C/C-SDSP-01.S",
    "rv64i_m/C/C-SLLI-01.S",
    "rv64i_m/C/C-SRAI-01.S",
    "rv64i_m/C/C-SRLI-01.S",
    "rv64i_m/C/C-SUB-01.S",
    "rv64i_m/C/C-SUBW-01.S",
    "rv64i_m/C/C-SW-01.S",
    "rv64i_m/C/C-SWSP-01.S",
    "rv64i_m/C/C-XOR-01.S",
    "rv64i_m/C/I-C-EBREAK-01.S",
    "rv64i_m/C/I-C-NOP-01.S"
  };

  string imperas64iNOc[] = {
    `IMPERASTEST,
    "rv64i_m/I/I-MISALIGN_JMP-01.S"
  };

  string imperas64i[] = '{
    `IMPERASTEST,
    "rv64i_m/I/I-DELAY_SLOTS-01.S",
    "rv64i_m/I/ADD-01.S",
    "rv64i_m/I/ADDI-01.S",
    "rv64i_m/I/ADDIW-01.S",
    "rv64i_m/I/ADDW-01.S",
    "rv64i_m/I/AND-01.S",
    "rv64i_m/I/ANDI-01.S",
    "rv64i_m/I/AUIPC-01.S",
    "rv64i_m/I/BEQ-01.S",
    "rv64i_m/I/BGE-01.S",
    "rv64i_m/I/BGEU-01.S",
    "rv64i_m/I/BLT-01.S",
    "rv64i_m/I/BLTU-01.S",
    "rv64i_m/I/BNE-01.S",
    "rv64i_m/I/I-DELAY_SLOTS-01.S",
    "rv64i_m/I/I-EBREAK-01.S",
    "rv64i_m/I/I-ECALL-01.S",
    "rv64i_m/I/I-ENDIANESS-01.S",
    "rv64i_m/I/I-IO-01.S",
//    "rv64i_m/I/I-MISALIGN_JMP-01.S",
    "rv64i_m/I/I-MISALIGN_LDST-01.S",
    "rv64i_m/I/I-NOP-01.S",
    "rv64i_m/I/I-RF_size-01.S",
    "rv64i_m/I/I-RF_width-01.S",
    "rv64i_m/I/I-RF_x0-01.S",
    "rv64i_m/I/JAL-01.S",
    "rv64i_m/I/JALR-01.S",
    "rv64i_m/I/LB-01.S",
    "rv64i_m/I/LBU-01.S",
    "rv64i_m/I/LD-01.S",
    "rv64i_m/I/LH-01.S",
    "rv64i_m/I/LHU-01.S",
    "rv64i_m/I/LUI-01.S",
    "rv64i_m/I/LW-01.S",
    "rv64i_m/I/LWU-01.S",
    "rv64i_m/I/OR-01.S",
    "rv64i_m/I/ORI-01.S",
    "rv64i_m/I/SB-01.S",
    "rv64i_m/I/SD-01.S",
    "rv64i_m/I/SH-01.S",
    "rv64i_m/I/SLL-01.S",
    "rv64i_m/I/SLLI-01.S",
    "rv64i_m/I/SLLIW-01.S",
    "rv64i_m/I/SLLW-01.S",
    "rv64i_m/I/SLT-01.S",
    "rv64i_m/I/SLTI-01.S",
    "rv64i_m/I/SLTIU-01.S",
    "rv64i_m/I/SLTU-01.S",
    "rv64i_m/I/SRA-01.S",
    "rv64i_m/I/SRAI-01.S",
    "rv64i_m/I/SRAIW-01.S",
    "rv64i_m/I/SRAW-01.S",
    "rv64i_m/I/SRL-01.S",
    "rv64i_m/I/SRLI-01.S",
    "rv64i_m/I/SRLIW-01.S",
    "rv64i_m/I/SRLW-01.S",
    "rv64i_m/I/SUB-01.S",
    "rv64i_m/I/SUBW-01.S",
    "rv64i_m/I/SW-01.S",
    "rv64i_m/I/XOR-01.S",
    "rv64i_m/I/XORI-01.S"
  };

  string imperas32m[] = '{
    `IMPERASTEST,
    "rv32i_m/M/DIV-01.S",
    "rv32i_m/M/DIVU-01.S",
    "rv32i_m/M/MUL-01.S",
    "rv32i_m/M/MULH-01.S",
    "rv32i_m/M/MULHSU-01.S",
    "rv32i_m/M/MULHU-01.S",
    "rv32i_m/M/REM-01.S",
    "rv32i_m/M/REMU-01.S"
  };

  string imperas32c[] = '{
    `IMPERASTEST,
    "rv32i_m/C/C-ADD-01.S",
    "rv32i_m/C/C-ADDI-01.S",
    "rv32i_m/C/C-ADDI16SP-01.S",
    "rv32i_m/C/C-ADDI4SPN-01.S",
    "rv32i_m/C/C-AND-01.S",
    "rv32i_m/C/C-ANDI-01.S",
    "rv32i_m/C/C-BEQZ-01.S",
    "rv32i_m/C/C-BNEZ-01.S",
    "rv32i_m/C/C-J-01.S",
    "rv32i_m/C/C-JAL-01.S",
    "rv32i_m/C/C-JALR-01.S",
    "rv32i_m/C/C-JR-01.S",
    "rv32i_m/C/C-LI-01.S",
    "rv32i_m/C/C-LUI-01.S",
    "rv32i_m/C/C-LW-01.S",
    "rv32i_m/C/C-LWSP-01.S",
    "rv32i_m/C/C-MV-01.S",
    "rv32i_m/C/C-OR-01.S",
    "rv32i_m/C/C-SLLI-01.S",
    "rv32i_m/C/C-SRAI-01.S",
    "rv32i_m/C/C-SRLI-01.S",
    "rv32i_m/C/C-SUB-01.S",
    "rv32i_m/C/C-SW-01.S",
    "rv32i_m/C/C-SWSP-01.S",
    "rv32i_m/C/C-XOR-01.S",
    "rv32i_m/C/I-C-EBREAK-01.S",
    "rv32i_m/C/I-C-NOP-01.S"
  };

  string imperas32iNOc[] = {
    `IMPERASTEST,
    "rv32i_m/I/I-MISALIGN_JMP-01.S"
  };

  string imperas32i[] = {
    `IMPERASTEST,
    "rv32i_m/I/ADD-01.S",
    "rv32i_m/I/ADDI-01.S",
    "rv32i_m/I/AND-01.S",
    "rv32i_m/I/ANDI-01.S",
    "rv32i_m/I/AUIPC-01.S",
    "rv32i_m/I/BEQ-01.S",
    "rv32i_m/I/BGE-01.S",
    "rv32i_m/I/BGEU-01.S",
    "rv32i_m/I/BLT-01.S",
    "rv32i_m/I/BLTU-01.S",
    "rv32i_m/I/BNE-01.S",
    "rv32i_m/I/I-DELAY_SLOTS-01.S",
    "rv32i_m/I/I-EBREAK-01.S",
    "rv32i_m/I/I-ECALL-01.S",
    "rv32i_m/I/I-ENDIANESS-01.S",
    "rv32i_m/I/I-IO-01.S",
//    "rv32i_m/I/I-MISALIGN_JMP-01.S",
    "rv32i_m/I/I-MISALIGN_LDST-01.S",
    "rv32i_m/I/I-NOP-01.S",
    "rv32i_m/I/I-RF_size-01.S",
    "rv32i_m/I/I-RF_width-01.S",
    "rv32i_m/I/I-RF_x0-01.S",
    "rv32i_m/I/JAL-01.S",
    "rv32i_m/I/JALR-01.S",
    "rv32i_m/I/LB-01.S",
    "rv32i_m/I/LBU-01.S",
    "rv32i_m/I/LH-01.S",
    "rv32i_m/I/LHU-01.S",
    "rv32i_m/I/LUI-01.S",
    "rv32i_m/I/LW-01.S",
    "rv32i_m/I/OR-01.S",
    "rv32i_m/I/ORI-01.S",
    "rv32i_m/I/SB-01.S",
    "rv32i_m/I/SH-01.S",
    "rv32i_m/I/SLL-01.S",
    "rv32i_m/I/SLLI-01.S",
    "rv32i_m/I/SLT-01.S",
    "rv32i_m/I/SLTI-01.S",
    "rv32i_m/I/SLTIU-01.S",
    "rv32i_m/I/SLTU-01.S",
    "rv32i_m/I/SRA-01.S",
    "rv32i_m/I/SRAI-01.S",
    "rv32i_m/I/SRL-01.S",
    "rv32i_m/I/SRLI-01.S",
    "rv32i_m/I/SUB-01.S",
    "rv32i_m/I/SW-01.S",
    "rv32i_m/I/XOR-01.S",
    "rv32i_m/I/XORI-01.S"   
  };


  string wally64a[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/src/WALLY-amo-01.S",
    "rv64i_m/privilege/src/WALLY-lrsc-01.S"
  };

  string wally32a[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/src/WALLY-amo-01.S",
    "rv32i_m/privilege/src/WALLY-lrsc-01.S"
    };

  string arch64priv[] = '{
    `RISCVARCHTEST,
    "rv64i_m/privilege/src/ebreak.S",
    "rv64i_m/privilege/src/ecall.S",
//    "rv64i_m/privilege/src/misalign1-jalr-01.S",
    "rv64i_m/privilege/src/misalign2-jalr-01.S",
    "rv64i_m/privilege/src/misalign-beq-01.S",
    "rv64i_m/privilege/src/misalign-bge-01.S",
    "rv64i_m/privilege/src/misalign-bgeu-01.S",
    "rv64i_m/privilege/src/misalign-blt-01.S",
    "rv64i_m/privilege/src/misalign-bltu-01.S",
    "rv64i_m/privilege/src/misalign-bne-01.S",
    "rv64i_m/privilege/src/misalign-jal-01.S",
    "rv64i_m/privilege/src/misalign-ld-01.S",
    "rv64i_m/privilege/src/misalign-lh-01.S",
    "rv64i_m/privilege/src/misalign-lhu-01.S",
    "rv64i_m/privilege/src/misalign-lw-01.S",
    "rv64i_m/privilege/src/misalign-lwu-01.S",
    "rv64i_m/privilege/src/misalign-sd-01.S",
    "rv64i_m/privilege/src/misalign-sh-01.S",
    "rv64i_m/privilege/src/misalign-sw-01.S"
    };

  string arch64zi[] = '{
    `RISCVARCHTEST,
    "rv64i_m/Zifencei/src/Fencei.S"
    };

  string arch32zi[] = '{
    `RISCVARCHTEST,
    "rv32i_m/Zifencei/src/Fencei.S"
    };

  string arch32zba[] = '{
    `RISCVARCHTEST,
    "rv32i_m/B/src/sh1add-01.S",
    "rv32i_m/B/src/sh2add-01.S",
    "rv32i_m/B/src/sh3add-01.S"
  };

  string arch32zbb[] = '{
    `RISCVARCHTEST,
    "rv32i_m/B/src/max-01.S",
    "rv32i_m/B/src/maxu-01.S",
    "rv32i_m/B/src/min-01.S",
    "rv32i_m/B/src/minu-01.S",
    "rv32i_m/B/src/orcb_32-01.S",
    "rv32i_m/B/src/rev8_32-01.S",
    "rv32i_m/B/src/andn-01.S",
    "rv32i_m/B/src/orn-01.S",
    "rv32i_m/B/src/xnor-01.S",
    "rv32i_m/B/src/zext.h_32-01.S",
    "rv32i_m/B/src/sext.b-01.S",
    "rv32i_m/B/src/sext.h-01.S",
    "rv32i_m/B/src/clz-01.S",
    "rv32i_m/B/src/cpop-01.S",
    "rv32i_m/B/src/ctz-01.S",
    "rv32i_m/B/src/ror-01.S",
    "rv32i_m/B/src/rori-01.S",
    "rv32i_m/B/src/rol-01.S"
  };

  string arch32zbc[] = '{
    `RISCVARCHTEST,
    "rv32i_m/B/src/clmul-01.S",
    "rv32i_m/B/src/clmulh-01.S",
    "rv32i_m/B/src/clmulr-01.S"
  };

  string arch32zbs[] = '{
    `RISCVARCHTEST,
    "rv32i_m/B/src/bclr-01.S",
    "rv32i_m/B/src/bclri-01.S",
    "rv32i_m/B/src/bext-01.S",
    "rv32i_m/B/src/bexti-01.S",
    "rv32i_m/B/src/binv-01.S",
    "rv32i_m/B/src/binvi-01.S",
    "rv32i_m/B/src/bset-01.S",
    "rv32i_m/B/src/bseti-01.S"
  };

  string arch32b[] = '{
    `RISCVARCHTEST,
    "rv32i_m/B/src/clmul-01.S",
    "rv32i_m/B/src/clmulh-01.S",
    "rv32i_m/B/src/clmulr-01.S",
    "rv32i_m/B/src/bclr-01.S",
    "rv32i_m/B/src/bclri-01.S",
    "rv32i_m/B/src/bext-01.S",
    "rv32i_m/B/src/bexti-01.S",
    "rv32i_m/B/src/binv-01.S",
    "rv32i_m/B/src/binvi-01.S",
    "rv32i_m/B/src/bset-01.S",
    "rv32i_m/B/src/bseti-01.S",
    "rv32i_m/B/src/max-01.S",
    "rv32i_m/B/src/maxu-01.S",
    "rv32i_m/B/src/min-01.S",
    "rv32i_m/B/src/minu-01.S",
    "rv32i_m/B/src/orcb_32-01.S",
    "rv32i_m/B/src/rev8_32-01.S",
    "rv32i_m/B/src/andn-01.S",
    "rv32i_m/B/src/orn-01.S",
    "rv32i_m/B/src/xnor-01.S",
    "rv32i_m/B/src/zext.h_32-01.S",
    "rv32i_m/B/src/sext.b-01.S",
    "rv32i_m/B/src/sext.h-01.S",
    "rv32i_m/B/src/clz-01.S",
    "rv32i_m/B/src/cpop-01.S",
    "rv32i_m/B/src/ctz-01.S",
    "rv32i_m/B/src/ror-01.S",
    "rv32i_m/B/src/rori-01.S",
    "rv32i_m/B/src/rol-01.S",
    "rv32i_m/B/src/sh1add-01.S",
    "rv32i_m/B/src/sh2add-01.S",
    "rv32i_m/B/src/sh3add-01.S",
    "rv32i_m/I/src/add-01.S",
    "rv32i_m/I/src/addi-01.S",
    "rv32i_m/I/src/and-01.S",
    "rv32i_m/I/src/andi-01.S",
    "rv32i_m/I/src/auipc-01.S",
    "rv32i_m/I/src/beq-01.S",
    "rv32i_m/I/src/bge-01.S",
    "rv32i_m/I/src/bgeu-01.S",
    "rv32i_m/I/src/blt-01.S",
    "rv32i_m/I/src/bltu-01.S",
    "rv32i_m/I/src/bne-01.S",
    "rv32i_m/I/src/fence-01.S",
    "rv32i_m/I/src/jal-01.S",
    "rv32i_m/I/src/jalr-01.S",
    "rv32i_m/I/src/lb-align-01.S",
    "rv32i_m/I/src/lbu-align-01.S",
    "rv32i_m/I/src/lh-align-01.S",
    "rv32i_m/I/src/lhu-align-01.S",
    "rv32i_m/I/src/lui-01.S",
    "rv32i_m/I/src/lw-align-01.S",
    "rv32i_m/I/src/or-01.S",
    "rv32i_m/I/src/ori-01.S",
    "rv32i_m/I/src/sb-align-01.S",
    "rv32i_m/I/src/sh-align-01.S",
    "rv32i_m/I/src/sll-01.S",
    "rv32i_m/I/src/slli-01.S",
    "rv32i_m/I/src/slt-01.S",
    "rv32i_m/I/src/slti-01.S",
    "rv32i_m/I/src/sltiu-01.S",
    "rv32i_m/I/src/sltu-01.S",
    "rv32i_m/I/src/sra-01.S",
    "rv32i_m/I/src/srai-01.S",
    "rv32i_m/I/src/srl-01.S",
    "rv32i_m/I/src/srli-01.S",
    "rv32i_m/I/src/sub-01.S",
    "rv32i_m/I/src/sw-align-01.S",
    "rv32i_m/I/src/xor-01.S",
    "rv32i_m/I/src/xori-01.S"
};

  string arch64m[] = '{
    `RISCVARCHTEST,
    "rv64i_m/M/src/div-01.S",
    "rv64i_m/M/src/divu-01.S",
    "rv64i_m/M/src/divuw-01.S",
    "rv64i_m/M/src/divw-01.S",
    "rv64i_m/M/src/mul-01.S",
    "rv64i_m/M/src/mulh-01.S",
    "rv64i_m/M/src/mulhsu-01.S",
    "rv64i_m/M/src/mulhu-01.S",
    "rv64i_m/M/src/mulw-01.S",
    "rv64i_m/M/src/rem-01.S",
    "rv64i_m/M/src/remu-01.S",
    "rv64i_m/M/src/remuw-01.S",
    "rv64i_m/M/src/remw-01.S"
   };

  string arch64c[] = '{
    `RISCVARCHTEST,
    "rv64i_m/C/src/cadd-01.S",
    "rv64i_m/C/src/caddi-01.S",
    "rv64i_m/C/src/caddi16sp-01.S",
    "rv64i_m/C/src/caddi4spn-01.S",
    "rv64i_m/C/src/caddiw-01.S",
    "rv64i_m/C/src/caddw-01.S",
    "rv64i_m/C/src/cand-01.S",
    "rv64i_m/C/src/candi-01.S",
    "rv64i_m/C/src/cbeqz-01.S",
    "rv64i_m/C/src/cbnez-01.S",
    "rv64i_m/C/src/cj-01.S",
    "rv64i_m/C/src/cjalr-01.S",
    "rv64i_m/C/src/cjr-01.S",
    "rv64i_m/C/src/cld-01.S",
    "rv64i_m/C/src/cldsp-01.S",
    "rv64i_m/C/src/cli-01.S",
    "rv64i_m/C/src/clui-01.S",
    "rv64i_m/C/src/clw-01.S",
    "rv64i_m/C/src/clwsp-01.S",
    "rv64i_m/C/src/cmv-01.S",
    "rv64i_m/C/src/cnop-01.S",
    "rv64i_m/C/src/cor-01.S",
    "rv64i_m/C/src/csd-01.S",
    "rv64i_m/C/src/csdsp-01.S",
    "rv64i_m/C/src/cslli-01.S",
    "rv64i_m/C/src/csrai-01.S",
    "rv64i_m/C/src/csrli-01.S",
    "rv64i_m/C/src/csub-01.S",
    "rv64i_m/C/src/csubw-01.S",
    "rv64i_m/C/src/csw-01.S",
    "rv64i_m/C/src/cswsp-01.S",
    "rv64i_m/C/src/cxor-01.S"
  };

  string arch64cpriv[] = '{
//    `RISCVARCHTEST,
    "rv64i_m/C/src/cebreak-01.S"
  };

  string arch64i[] = '{
    `RISCVARCHTEST,
    "rv64i_m/I/src/add-01.S",
    "rv64i_m/I/src/addi-01.S",
    "rv64i_m/I/src/addiw-01.S",
    "rv64i_m/I/src/addw-01.S",
    "rv64i_m/I/src/and-01.S",
    "rv64i_m/I/src/andi-01.S",
    "rv64i_m/I/src/auipc-01.S",
    "rv64i_m/I/src/beq-01.S",
    "rv64i_m/I/src/bge-01.S",
    "rv64i_m/I/src/bgeu-01.S",
    "rv64i_m/I/src/blt-01.S",
    "rv64i_m/I/src/bltu-01.S",
    "rv64i_m/I/src/bne-01.S",
    "rv64i_m/I/src/fence-01.S",
    "rv64i_m/I/src/jal-01.S",
    "rv64i_m/I/src/jalr-01.S",
    "rv64i_m/I/src/lb-align-01.S",
    "rv64i_m/I/src/lbu-align-01.S",
    "rv64i_m/I/src/ld-align-01.S",
    "rv64i_m/I/src/lh-align-01.S",
    "rv64i_m/I/src/lhu-align-01.S",
    "rv64i_m/I/src/lui-01.S",
    "rv64i_m/I/src/lw-align-01.S",
    "rv64i_m/I/src/lwu-align-01.S",
    "rv64i_m/I/src/or-01.S",
    "rv64i_m/I/src/ori-01.S",
    "rv64i_m/I/src/sb-align-01.S",
    "rv64i_m/I/src/sd-align-01.S",
    "rv64i_m/I/src/sh-align-01.S",
    "rv64i_m/I/src/sll-01.S",
    "rv64i_m/I/src/slli-01.S",
    "rv64i_m/I/src/slliw-01.S",
    "rv64i_m/I/src/sllw-01.S",
    "rv64i_m/I/src/slt-01.S",
    "rv64i_m/I/src/slti-01.S",
    "rv64i_m/I/src/sltiu-01.S",
    "rv64i_m/I/src/sltu-01.S",
    "rv64i_m/I/src/sra-01.S",
    "rv64i_m/I/src/srai-01.S",
    "rv64i_m/I/src/sraiw-01.S",
    "rv64i_m/I/src/sraw-01.S",
    "rv64i_m/I/src/srl-01.S",
    "rv64i_m/I/src/srli-01.S",
    "rv64i_m/I/src/srliw-01.S",
    "rv64i_m/I/src/srlw-01.S",
    "rv64i_m/I/src/sub-01.S",
    "rv64i_m/I/src/subw-01.S",
    "rv64i_m/I/src/sw-align-01.S",
    "rv64i_m/I/src/xor-01.S",
    "rv64i_m/I/src/xori-01.S"
  };

  string arch64f[] = '{
    `RISCVARCHTEST,
    "rv64i_m/F/src/fadd_b10-01.S",
    "rv64i_m/F/src/fadd_b1-01.S",
    "rv64i_m/F/src/fadd_b11-01.S",
    "rv64i_m/F/src/fadd_b12-01.S",
    "rv64i_m/F/src/fadd_b13-01.S",
    "rv64i_m/F/src/fadd_b2-01.S",
    "rv64i_m/F/src/fadd_b3-01.S",
    "rv64i_m/F/src/fadd_b4-01.S",
    "rv64i_m/F/src/fadd_b5-01.S",
    "rv64i_m/F/src/fadd_b7-01.S",
    "rv64i_m/F/src/fadd_b8-01.S",
    "rv64i_m/F/src/fclass_b1-01.S",
    "rv64i_m/F/src/fcvt.s.w_b25-01.S",
    "rv64i_m/F/src/fcvt.s.w_b26-01.S",
    "rv64i_m/F/src/fcvt.s.wu_b25-01.S",
    "rv64i_m/F/src/fcvt.s.wu_b26-01.S",
    "rv64i_m/F/src/fcvt.w.s_b1-01.S",
    "rv64i_m/F/src/fcvt.w.s_b22-01.S",
    "rv64i_m/F/src/fcvt.w.s_b23-01.S",
    "rv64i_m/F/src/fcvt.w.s_b24-01.S",
    "rv64i_m/F/src/fcvt.w.s_b27-01.S",
    "rv64i_m/F/src/fcvt.w.s_b28-01.S",
    "rv64i_m/F/src/fcvt.w.s_b29-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b1-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b22-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b23-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b24-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b27-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b28-01.S",
    "rv64i_m/F/src/fcvt.wu.s_b29-01.S",
    "rv64i_m/F/src/fdiv_b1-01.S",
    "rv64i_m/F/src/fdiv_b20-01.S",
    "rv64i_m/F/src/fdiv_b2-01.S",
    "rv64i_m/F/src/fdiv_b21-01.S",
    "rv64i_m/F/src/fdiv_b3-01.S",
    "rv64i_m/F/src/fdiv_b4-01.S",
    "rv64i_m/F/src/fdiv_b5-01.S",
    "rv64i_m/F/src/fdiv_b6-01.S",
    "rv64i_m/F/src/fdiv_b7-01.S",
    "rv64i_m/F/src/fdiv_b8-01.S",
    "rv64i_m/F/src/fdiv_b9-01.S",
    "rv64i_m/F/src/feq_b1-01.S",
    "rv64i_m/F/src/feq_b19-01.S",
    "rv64i_m/F/src/fle_b1-01.S",
    "rv64i_m/F/src/fle_b19-01.S",
    "rv64i_m/F/src/flt_b1-01.S",
    "rv64i_m/F/src/flt_b19-01.S",
    "rv64i_m/F/src/flw-align-01.S",
    "rv64i_m/F/src/fmadd_b1-01.S",
    "rv64i_m/F/src/fmadd_b14-01.S",
    //"rv64i_m/F/src/fmadd_b15-01.S",
    "rv64i_m/F/src/fmadd_b16-01.S",
    "rv64i_m/F/src/fmadd_b17-01.S",
    "rv64i_m/F/src/fmadd_b18-01.S",
    "rv64i_m/F/src/fmadd_b2-01.S",
    "rv64i_m/F/src/fmadd_b3-01.S",
    "rv64i_m/F/src/fmadd_b4-01.S",
    "rv64i_m/F/src/fmadd_b5-01.S",
    "rv64i_m/F/src/fmadd_b6-01.S",
    "rv64i_m/F/src/fmadd_b7-01.S",
    "rv64i_m/F/src/fmadd_b8-01.S",
    "rv64i_m/F/src/fmax_b1-01.S",
    "rv64i_m/F/src/fmax_b19-01.S",
    "rv64i_m/F/src/fmin_b1-01.S",
    "rv64i_m/F/src/fmin_b19-01.S",
    "rv64i_m/F/src/fmsub_b1-01.S",
    "rv64i_m/F/src/fmsub_b14-01.S",
    "rv64i_m/F/src/fmsub_b15-01.S",
    "rv64i_m/F/src/fmsub_b16-01.S",
    "rv64i_m/F/src/fmsub_b17-01.S",
    "rv64i_m/F/src/fmsub_b18-01.S",
    "rv64i_m/F/src/fmsub_b2-01.S",
    "rv64i_m/F/src/fmsub_b3-01.S",
    "rv64i_m/F/src/fmsub_b4-01.S",
    "rv64i_m/F/src/fmsub_b5-01.S",
    "rv64i_m/F/src/fmsub_b6-01.S",
    "rv64i_m/F/src/fmsub_b7-01.S",
    "rv64i_m/F/src/fmsub_b8-01.S",
    "rv64i_m/F/src/fmul_b1-01.S",
    "rv64i_m/F/src/fmul_b2-01.S",
    "rv64i_m/F/src/fmul_b3-01.S",
    "rv64i_m/F/src/fmul_b4-01.S",
    "rv64i_m/F/src/fmul_b5-01.S",
    "rv64i_m/F/src/fmul_b6-01.S",
    "rv64i_m/F/src/fmul_b7-01.S",
    "rv64i_m/F/src/fmul_b8-01.S",
    "rv64i_m/F/src/fmul_b9-01.S",
    "rv64i_m/F/src/fmv.w.x_b25-01.S",
    "rv64i_m/F/src/fmv.w.x_b26-01.S",
    "rv64i_m/F/src/fmv.x.w_b1-01.S",
    "rv64i_m/F/src/fmv.x.w_b22-01.S",
    "rv64i_m/F/src/fmv.x.w_b23-01.S",
    "rv64i_m/F/src/fmv.x.w_b24-01.S",
    "rv64i_m/F/src/fmv.x.w_b27-01.S",
    "rv64i_m/F/src/fmv.x.w_b28-01.S",
    "rv64i_m/F/src/fmv.x.w_b29-01.S",
    "rv64i_m/F/src/fnmadd_b1-01.S",
    "rv64i_m/F/src/fnmadd_b14-01.S",
    // "rv64i_m/F/src/fnmadd_b15-01.S",
    "rv64i_m/F/src/fnmadd_b16-01.S",
    "rv64i_m/F/src/fnmadd_b17-01.S",
    "rv64i_m/F/src/fnmadd_b18-01.S",
    "rv64i_m/F/src/fnmadd_b2-01.S",
    "rv64i_m/F/src/fnmadd_b3-01.S",
    "rv64i_m/F/src/fnmadd_b4-01.S",
    "rv64i_m/F/src/fnmadd_b5-01.S",
    "rv64i_m/F/src/fnmadd_b6-01.S",
    "rv64i_m/F/src/fnmadd_b7-01.S",
    "rv64i_m/F/src/fnmadd_b8-01.S",
    "rv64i_m/F/src/fnmsub_b1-01.S",
    "rv64i_m/F/src/fnmsub_b14-01.S",
    // "rv64i_m/F/src/fnmsub_b15-01.S",
    "rv64i_m/F/src/fnmsub_b16-01.S",
    "rv64i_m/F/src/fnmsub_b17-01.S",
    "rv64i_m/F/src/fnmsub_b18-01.S",
    "rv64i_m/F/src/fnmsub_b2-01.S",
    "rv64i_m/F/src/fnmsub_b3-01.S",
    "rv64i_m/F/src/fnmsub_b4-01.S",
    "rv64i_m/F/src/fnmsub_b5-01.S",
    "rv64i_m/F/src/fnmsub_b6-01.S",
    "rv64i_m/F/src/fnmsub_b7-01.S",
    "rv64i_m/F/src/fnmsub_b8-01.S",
    "rv64i_m/F/src/fsgnj_b1-01.S",
    "rv64i_m/F/src/fsgnjn_b1-01.S",
    "rv64i_m/F/src/fsgnjx_b1-01.S",
    "rv64i_m/F/src/fsqrt_b1-01.S",
    "rv64i_m/F/src/fsqrt_b20-01.S",
    "rv64i_m/F/src/fsqrt_b2-01.S",
    "rv64i_m/F/src/fsqrt_b3-01.S",
    "rv64i_m/F/src/fsqrt_b4-01.S",
    "rv64i_m/F/src/fsqrt_b5-01.S",
    "rv64i_m/F/src/fsqrt_b7-01.S",
    "rv64i_m/F/src/fsqrt_b8-01.S",
    "rv64i_m/F/src/fsqrt_b9-01.S",
    "rv64i_m/F/src/fsub_b10-01.S",
    "rv64i_m/F/src/fsub_b1-01.S",
    "rv64i_m/F/src/fsub_b11-01.S",
    "rv64i_m/F/src/fsub_b12-01.S",
    "rv64i_m/F/src/fsub_b13-01.S",
    "rv64i_m/F/src/fsub_b2-01.S",
    "rv64i_m/F/src/fsub_b3-01.S",
    "rv64i_m/F/src/fsub_b4-01.S",
    "rv64i_m/F/src/fsub_b5-01.S",
    "rv64i_m/F/src/fsub_b7-01.S",
    "rv64i_m/F/src/fsub_b8-01.S",
    "rv64i_m/F/src/fsw-align-01.S"
    };


  string arch64d[] = '{
    `RISCVARCHTEST,
    "rv64i_m/D/src/fadd.d_b10-01.S",
    "rv64i_m/D/src/fadd.d_b1-01.S",
    "rv64i_m/D/src/fadd.d_b11-01.S",
    "rv64i_m/D/src/fadd.d_b12-01.S",
    "rv64i_m/D/src/fadd.d_b13-01.S",
    "rv64i_m/D/src/fadd.d_b2-01.S",
    "rv64i_m/D/src/fadd.d_b3-01.S",
    "rv64i_m/D/src/fadd.d_b4-01.S",
    "rv64i_m/D/src/fadd.d_b5-01.S",
    "rv64i_m/D/src/fadd.d_b7-01.S",
    "rv64i_m/D/src/fadd.d_b8-01.S",
    "rv64i_m/D/src/fclass.d_b1-01.S",
    "rv64i_m/D/src/fcvt.d.l_b25-01.S",
    "rv64i_m/D/src/fcvt.d.l_b26-01.S",
    "rv64i_m/D/src/fcvt.d.lu_b25-01.S",
    "rv64i_m/D/src/fcvt.d.lu_b26-01.S",
    "rv64i_m/D/src/fcvt.d.s_b1-01.S",
    "rv64i_m/D/src/fcvt.d.s_b22-01.S",
    "rv64i_m/D/src/fcvt.d.s_b23-01.S",
    "rv64i_m/D/src/fcvt.d.s_b24-01.S",
    "rv64i_m/D/src/fcvt.d.s_b27-01.S",
    "rv64i_m/D/src/fcvt.d.s_b28-01.S",
    "rv64i_m/D/src/fcvt.d.s_b29-01.S",
    "rv64i_m/D/src/fcvt.d.w_b25-01.S",
    "rv64i_m/D/src/fcvt.d.w_b26-01.S",
    "rv64i_m/D/src/fcvt.d.wu_b25-01.S",
    "rv64i_m/D/src/fcvt.d.wu_b26-01.S",
    "rv64i_m/D/src/fcvt.l.d_b1-01.S",
    "rv64i_m/D/src/fcvt.l.d_b22-01.S",
    "rv64i_m/D/src/fcvt.l.d_b23-01.S",
    "rv64i_m/D/src/fcvt.l.d_b24-01.S",
    "rv64i_m/D/src/fcvt.l.d_b27-01.S",
    "rv64i_m/D/src/fcvt.l.d_b28-01.S",
    "rv64i_m/D/src/fcvt.l.d_b29-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b1-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b22-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b23-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b24-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b27-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b28-01.S",
    "rv64i_m/D/src/fcvt.lu.d_b29-01.S",
    "rv64i_m/D/src/fcvt.s.d_b1-01.S",
    "rv64i_m/D/src/fcvt.s.d_b22-01.S",
    "rv64i_m/D/src/fcvt.s.d_b23-01.S",
    "rv64i_m/D/src/fcvt.s.d_b24-01.S",
    "rv64i_m/D/src/fcvt.s.d_b27-01.S",
    "rv64i_m/D/src/fcvt.s.d_b28-01.S",
    "rv64i_m/D/src/fcvt.s.d_b29-01.S",
    "rv64i_m/D/src/fcvt.w.d_b1-01.S",
    "rv64i_m/D/src/fcvt.w.d_b22-01.S",
    "rv64i_m/D/src/fcvt.w.d_b23-01.S",
    "rv64i_m/D/src/fcvt.w.d_b24-01.S",
    "rv64i_m/D/src/fcvt.w.d_b27-01.S",
    "rv64i_m/D/src/fcvt.w.d_b28-01.S",
    "rv64i_m/D/src/fcvt.w.d_b29-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b1-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b22-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b23-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b24-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b27-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b28-01.S",
    "rv64i_m/D/src/fcvt.wu.d_b29-01.S",
    "rv64i_m/D/src/fdiv.d_b1-01.S",
    "rv64i_m/D/src/fdiv.d_b20-01.S",
    "rv64i_m/D/src/fdiv.d_b2-01.S",
    "rv64i_m/D/src/fdiv.d_b21-01.S",
    "rv64i_m/D/src/fdiv.d_b3-01.S",
    "rv64i_m/D/src/fdiv.d_b4-01.S",
    "rv64i_m/D/src/fdiv.d_b5-01.S",
    "rv64i_m/D/src/fdiv.d_b6-01.S",
    "rv64i_m/D/src/fdiv.d_b7-01.S",
    "rv64i_m/D/src/fdiv.d_b8-01.S",
    "rv64i_m/D/src/fdiv.d_b9-01.S",
    "rv64i_m/D/src/feq.d_b1-01.S",
    "rv64i_m/D/src/feq.d_b19-01.S",
    "rv64i_m/D/src/fle.d_b1-01.S",
    "rv64i_m/D/src/fle.d_b19-01.S",
    "rv64i_m/D/src/flt.d_b1-01.S",
    "rv64i_m/D/src/flt.d_b19-01.S",
    "rv64i_m/D/src/fld-align-01.S", 
    "rv64i_m/D/src/fsd-align-01.S", 
    "rv64i_m/D/src/fmadd.d_b14-01.S",
    "rv64i_m/D/src/fmadd.d_b16-01.S",
    "rv64i_m/D/src/fmadd.d_b17-01.S",
    "rv64i_m/D/src/fmadd.d_b18-01.S",
    "rv64i_m/D/src/fmadd.d_b2-01.S",
    "rv64i_m/D/src/fmadd.d_b3-01.S",
    "rv64i_m/D/src/fmadd.d_b4-01.S",
    "rv64i_m/D/src/fmadd.d_b5-01.S",
    "rv64i_m/D/src/fmadd.d_b6-01.S",
    "rv64i_m/D/src/fmadd.d_b7-01.S",
    "rv64i_m/D/src/fmadd.d_b8-01.S",
    "rv64i_m/D/src/fmax.d_b1-01.S",
    "rv64i_m/D/src/fmax.d_b19-01.S",
    "rv64i_m/D/src/fmin.d_b1-01.S",
    "rv64i_m/D/src/fmin.d_b19-01.S",
    "rv64i_m/D/src/fmsub.d_b14-01.S",
    "rv64i_m/D/src/fmsub.d_b16-01.S",
    "rv64i_m/D/src/fmsub.d_b17-01.S",
    "rv64i_m/D/src/fmsub.d_b18-01.S",
    "rv64i_m/D/src/fmsub.d_b2-01.S",
    "rv64i_m/D/src/fmsub.d_b3-01.S",
    "rv64i_m/D/src/fmsub.d_b4-01.S",
    "rv64i_m/D/src/fmsub.d_b5-01.S",
    "rv64i_m/D/src/fmsub.d_b6-01.S",
    "rv64i_m/D/src/fmsub.d_b7-01.S",
    "rv64i_m/D/src/fmsub.d_b8-01.S",
    "rv64i_m/D/src/fmul.d_b1-01.S",
    "rv64i_m/D/src/fmul.d_b2-01.S",
    "rv64i_m/D/src/fmul.d_b3-01.S",
    "rv64i_m/D/src/fmul.d_b4-01.S",
    "rv64i_m/D/src/fmul.d_b5-01.S",
    "rv64i_m/D/src/fmul.d_b6-01.S",
    "rv64i_m/D/src/fmul.d_b7-01.S",
    "rv64i_m/D/src/fmul.d_b8-01.S",
    "rv64i_m/D/src/fmul.d_b9-01.S",
    "rv64i_m/D/src/fmv.d.x_b25-01.S",
    "rv64i_m/D/src/fmv.d.x_b26-01.S",
    "rv64i_m/D/src/fmv.x.d_b1-01.S",
    "rv64i_m/D/src/fmv.x.d_b22-01.S",
    "rv64i_m/D/src/fmv.x.d_b23-01.S",
    "rv64i_m/D/src/fmv.x.d_b24-01.S",
    "rv64i_m/D/src/fmv.x.d_b27-01.S",
    "rv64i_m/D/src/fmv.x.d_b28-01.S",
    "rv64i_m/D/src/fmv.x.d_b29-01.S",
    "rv64i_m/D/src/fnmadd.d_b14-01.S",
    "rv64i_m/D/src/fnmadd.d_b16-01.S",
    "rv64i_m/D/src/fnmadd.d_b17-01.S",
    "rv64i_m/D/src/fnmadd.d_b18-01.S",
    "rv64i_m/D/src/fnmadd.d_b2-01.S",
    "rv64i_m/D/src/fnmadd.d_b3-01.S",
    "rv64i_m/D/src/fnmadd.d_b4-01.S",
    "rv64i_m/D/src/fnmadd.d_b5-01.S",
    "rv64i_m/D/src/fnmadd.d_b6-01.S",
    "rv64i_m/D/src/fnmadd.d_b7-01.S",
    "rv64i_m/D/src/fnmadd.d_b8-01.S",
    "rv64i_m/D/src/fnmsub.d_b14-01.S",
    "rv64i_m/D/src/fnmsub.d_b16-01.S",
    "rv64i_m/D/src/fnmsub.d_b17-01.S",
    "rv64i_m/D/src/fnmsub.d_b18-01.S",
    "rv64i_m/D/src/fnmsub.d_b2-01.S",
    "rv64i_m/D/src/fnmsub.d_b3-01.S",
    "rv64i_m/D/src/fnmsub.d_b4-01.S",
    "rv64i_m/D/src/fnmsub.d_b5-01.S",
    "rv64i_m/D/src/fnmsub.d_b6-01.S",
    "rv64i_m/D/src/fnmsub.d_b7-01.S",
    "rv64i_m/D/src/fnmsub.d_b8-01.S",
    "rv64i_m/D/src/fsgnj.d_b1-01.S",
    "rv64i_m/D/src/fsgnjn.d_b1-01.S",
    "rv64i_m/D/src/fsgnjx.d_b1-01.S",
    "rv64i_m/D/src/fsqrt.d_b1-01.S",
    "rv64i_m/D/src/fsqrt.d_b20-01.S",
    "rv64i_m/D/src/fsqrt.d_b2-01.S",
    "rv64i_m/D/src/fsqrt.d_b3-01.S",
    "rv64i_m/D/src/fsqrt.d_b4-01.S",
    "rv64i_m/D/src/fsqrt.d_b5-01.S",
    "rv64i_m/D/src/fsqrt.d_b7-01.S",
    "rv64i_m/D/src/fsqrt.d_b8-01.S",
    "rv64i_m/D/src/fsqrt.d_b9-01.S",
    "rv64i_m/D/src/fssub.d_b10-01.S",
    "rv64i_m/D/src/fssub.d_b1-01.S",
    "rv64i_m/D/src/fssub.d_b11-01.S",
    "rv64i_m/D/src/fssub.d_b12-01.S",
    "rv64i_m/D/src/fssub.d_b13-01.S",
    "rv64i_m/D/src/fssub.d_b2-01.S",
    "rv64i_m/D/src/fssub.d_b3-01.S",
    "rv64i_m/D/src/fssub.d_b4-01.S",
    "rv64i_m/D/src/fssub.d_b5-01.S",
    "rv64i_m/D/src/fssub.d_b7-01.S",
    "rv64i_m/D/src/fssub.d_b8-01.S"
};


string arch64b[] = '{
    `RISCVARCHTEST,
    "rv64i_m/B/src/max-01.S",
    "rv64i_m/B/src/maxu-01.S",
    "rv64i_m/B/src/min-01.S",
    "rv64i_m/B/src/minu-01.S",
    "rv64i_m/B/src/orcb_64-01.S",
    "rv64i_m/B/src/rev8-01.S",
    "rv64i_m/B/src/andn-01.S",
    "rv64i_m/B/src/orn-01.S",
    "rv64i_m/B/src/xnor-01.S",
    "rv64i_m/B/src/zext.h-01.S",
    "rv64i_m/B/src/sext.b-01.S",
    "rv64i_m/B/src/sext.h-01.S",
    "rv64i_m/B/src/clz-01.S",
    "rv64i_m/B/src/clzw-01.S",
    "rv64i_m/B/src/cpop-01.S",
    "rv64i_m/B/src/cpopw-01.S",
    "rv64i_m/B/src/ctz-01.S",
    "rv64i_m/B/src/ctzw-01.S",
    "rv64i_m/B/src/rolw-01.S",
    "rv64i_m/B/src/ror-01.S",
    "rv64i_m/B/src/rori-01.S",
    "rv64i_m/B/src/roriw-01.S",
    "rv64i_m/B/src/rorw-01.S",
    "rv64i_m/B/src/rol-01.S",
    "rv64i_m/B/src/slli.uw-01.S",
    "rv64i_m/B/src/add.uw-01.S",
    "rv64i_m/B/src/sh1add-01.S",
    "rv64i_m/B/src/sh2add-01.S",
    "rv64i_m/B/src/sh3add-01.S",
    "rv64i_m/B/src/sh1add.uw-01.S",
    "rv64i_m/B/src/sh2add.uw-01.S",
    "rv64i_m/B/src/sh3add.uw-01.S",
    "rv64i_m/I/src/add-01.S",
    "rv64i_m/I/src/addi-01.S",
    "rv64i_m/I/src/addiw-01.S",
    "rv64i_m/I/src/addw-01.S",
    "rv64i_m/I/src/and-01.S",
    "rv64i_m/I/src/andi-01.S",
    "rv64i_m/I/src/auipc-01.S",
    "rv64i_m/I/src/beq-01.S",
    "rv64i_m/I/src/bge-01.S",
    "rv64i_m/I/src/bgeu-01.S",
    "rv64i_m/I/src/blt-01.S",
    "rv64i_m/I/src/bltu-01.S",
    "rv64i_m/I/src/bne-01.S",
    "rv64i_m/I/src/fence-01.S",
    "rv64i_m/I/src/jal-01.S",
    "rv64i_m/I/src/jalr-01.S",
    "rv64i_m/I/src/lb-align-01.S",
    "rv64i_m/I/src/lbu-align-01.S",
    "rv64i_m/I/src/ld-align-01.S",
    "rv64i_m/I/src/lh-align-01.S",
    "rv64i_m/I/src/lhu-align-01.S",
    "rv64i_m/I/src/lui-01.S",
    "rv64i_m/I/src/lw-align-01.S",
    "rv64i_m/I/src/lwu-align-01.S",
    "rv64i_m/I/src/or-01.S",
    "rv64i_m/I/src/ori-01.S",
    "rv64i_m/I/src/sb-align-01.S",
    "rv64i_m/I/src/sd-align-01.S",
    "rv64i_m/I/src/sh-align-01.S",
    "rv64i_m/I/src/sll-01.S",
    "rv64i_m/I/src/slli-01.S",
    "rv64i_m/I/src/slliw-01.S",
    "rv64i_m/I/src/sllw-01.S",
    "rv64i_m/I/src/slt-01.S",
    "rv64i_m/I/src/slti-01.S",
    "rv64i_m/I/src/sltiu-01.S",
    "rv64i_m/I/src/sltu-01.S",
    "rv64i_m/I/src/sra-01.S",
    "rv64i_m/I/src/srai-01.S",
    "rv64i_m/I/src/sraiw-01.S",
    "rv64i_m/I/src/sraw-01.S",
    "rv64i_m/I/src/srl-01.S",
    "rv64i_m/I/src/srli-01.S",
    "rv64i_m/I/src/srliw-01.S",
    "rv64i_m/I/src/srlw-01.S",
    "rv64i_m/I/src/sub-01.S",
    "rv64i_m/I/src/subw-01.S",
    "rv64i_m/I/src/sw-align-01.S",
    "rv64i_m/I/src/xor-01.S",
    "rv64i_m/I/src/xori-01.S",
    "rv64i_m/B/src/clmul-01.S",
    "rv64i_m/B/src/clmulh-01.S",
    "rv64i_m/B/src/clmulr-01.S",
    "rv64i_m/B/src/bclr-01.S",
    "rv64i_m/B/src/bclri-01.S",
    "rv64i_m/B/src/bext-01.S",
    "rv64i_m/B/src/bexti-01.S",
    "rv64i_m/B/src/binv-01.S",
    "rv64i_m/B/src/binvi-01.S",
    "rv64i_m/B/src/bset-01.S",
    "rv64i_m/B/src/bseti-01.S"
};

  string arch64zba[] = '{
      `RISCVARCHTEST,
      "rv64i_m/B/src/slli.uw-01.S",
      "rv64i_m/B/src/add.uw-01.S",
      "rv64i_m/B/src/sh1add-01.S",
      "rv64i_m/B/src/sh2add-01.S",
      "rv64i_m/B/src/sh3add-01.S",
      "rv64i_m/B/src/sh1add.uw-01.S",
      "rv64i_m/B/src/sh2add.uw-01.S",
      "rv64i_m/B/src/sh3add.uw-01.S"
  };



string arch64zbb[] = '{
    `RISCVARCHTEST,
    "rv64i_m/B/src/max-01.S",
    "rv64i_m/B/src/maxu-01.S",
    "rv64i_m/B/src/min-01.S",
    "rv64i_m/B/src/minu-01.S",
    "rv64i_m/B/src/orcb_64-01.S",
    "rv64i_m/B/src/rev8-01.S",
    "rv64i_m/B/src/andn-01.S",
    "rv64i_m/B/src/orn-01.S",
    "rv64i_m/B/src/xnor-01.S",
    "rv64i_m/B/src/zext.h-01.S",
    "rv64i_m/B/src/sext.b-01.S",
    "rv64i_m/B/src/sext.h-01.S",
    "rv64i_m/B/src/clz-01.S",
    "rv64i_m/B/src/clzw-01.S",
    "rv64i_m/B/src/cpop-01.S",
    "rv64i_m/B/src/cpopw-01.S",
    "rv64i_m/B/src/ctz-01.S",
    "rv64i_m/B/src/ctzw-01.S",
    "rv64i_m/B/src/rolw-01.S",
    "rv64i_m/B/src/ror-01.S",
    "rv64i_m/B/src/rori-01.S",
    "rv64i_m/B/src/roriw-01.S",
    "rv64i_m/B/src/rorw-01.S",
    "rv64i_m/B/src/rol-01.S"
};

string arch64zbc[] = '{
    `RISCVARCHTEST,
    "rv64i_m/B/src/clmul-01.S",
    "rv64i_m/B/src/clmulh-01.S",
    "rv64i_m/B/src/clmulr-01.S"
};

string arch64zbs[] = '{
    `RISCVARCHTEST,
    "rv64i_m/B/src/bclr-01.S",
    "rv64i_m/B/src/bclri-01.S",
    "rv64i_m/B/src/bext-01.S",
    "rv64i_m/B/src/bexti-01.S",
    "rv64i_m/B/src/binv-01.S",
    "rv64i_m/B/src/binvi-01.S",
    "rv64i_m/B/src/bset-01.S",
    "rv64i_m/B/src/bseti-01.S"
};



    string arch32priv[] = '{
    `RISCVARCHTEST,
    "rv32i_m/privilege/src/ebreak.S",
    "rv32i_m/privilege/src/ecall.S",
//    "rv32i_m/privilege/src/misalign1-jalr-01.S",
    "rv32i_m/privilege/src/misalign2-jalr-01.S",
    "rv32i_m/privilege/src/misalign-beq-01.S",
    "rv32i_m/privilege/src/misalign-bge-01.S",
    "rv32i_m/privilege/src/misalign-bgeu-01.S",
    "rv32i_m/privilege/src/misalign-blt-01.S",
    "rv32i_m/privilege/src/misalign-bltu-01.S",
    "rv32i_m/privilege/src/misalign-bne-01.S",
    "rv32i_m/privilege/src/misalign-jal-01.S",
    "rv32i_m/privilege/src/misalign-lh-01.S",
    "rv32i_m/privilege/src/misalign-lhu-01.S",
    "rv32i_m/privilege/src/misalign-lw-01.S",
    "rv32i_m/privilege/src/misalign-sh-01.S",
    "rv32i_m/privilege/src/misalign-sw-01.S"
    };

  string arch32m[] = '{
    `RISCVARCHTEST,
    "rv32i_m/M/src/div-01.S",
    "rv32i_m/M/src/divu-01.S",
    "rv32i_m/M/src/rem-01.S",
    "rv32i_m/M/src/remu-01.S",
    "rv32i_m/M/src/mul-01.S",
    "rv32i_m/M/src/mulh-01.S",
    "rv32i_m/M/src/mulhsu-01.S",
    "rv32i_m/M/src/mulhu-01.S"
   };

  string arch32f[] = '{
    `RISCVARCHTEST,
    "rv32i_m/F/src/fdiv_b20-01.S",
    "rv32i_m/F/src/fadd_b10-01.S",
    "rv32i_m/F/src/fadd_b1-01.S",
    "rv32i_m/F/src/fadd_b11-01.S",
    "rv32i_m/F/src/fadd_b12-01.S",
    "rv32i_m/F/src/fadd_b13-01.S",
    "rv32i_m/F/src/fadd_b2-01.S",
    "rv32i_m/F/src/fadd_b3-01.S",
    "rv32i_m/F/src/fadd_b4-01.S",
    "rv32i_m/F/src/fadd_b5-01.S",
    "rv32i_m/F/src/fadd_b7-01.S",
    "rv32i_m/F/src/fadd_b8-01.S",
    "rv32i_m/F/src/fclass_b1-01.S",
    "rv32i_m/F/src/fcvt.s.w_b25-01.S",
    "rv32i_m/F/src/fcvt.s.w_b26-01.S",
    "rv32i_m/F/src/fcvt.s.wu_b25-01.S",
    "rv32i_m/F/src/fcvt.s.wu_b26-01.S",
    "rv32i_m/F/src/fcvt.w.s_b1-01.S",
    "rv32i_m/F/src/fcvt.w.s_b22-01.S",
    "rv32i_m/F/src/fcvt.w.s_b23-01.S",
    "rv32i_m/F/src/fcvt.w.s_b24-01.S",
    "rv32i_m/F/src/fcvt.w.s_b27-01.S",
    "rv32i_m/F/src/fcvt.w.s_b28-01.S",
    "rv32i_m/F/src/fcvt.w.s_b29-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b1-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b22-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b23-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b24-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b27-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b28-01.S",
    "rv32i_m/F/src/fcvt.wu.s_b29-01.S",
    "rv32i_m/F/src/fdiv_b20-01.S",
    "rv32i_m/F/src/fdiv_b1-01.S",
    "rv32i_m/F/src/fdiv_b2-01.S",
    "rv32i_m/F/src/fdiv_b21-01.S",
    "rv32i_m/F/src/fdiv_b3-01.S",
    "rv32i_m/F/src/fdiv_b4-01.S",
    "rv32i_m/F/src/fdiv_b5-01.S",
    "rv32i_m/F/src/fdiv_b6-01.S",
    "rv32i_m/F/src/fdiv_b7-01.S",
    "rv32i_m/F/src/fdiv_b8-01.S",
    "rv32i_m/F/src/fdiv_b9-01.S",
    "rv32i_m/F/src/feq_b1-01.S",
    "rv32i_m/F/src/feq_b19-01.S",
    "rv32i_m/F/src/fle_b1-01.S",
    "rv32i_m/F/src/fle_b19-01.S",
    "rv32i_m/F/src/flt_b1-01.S",
    "rv32i_m/F/src/flt_b19-01.S",
    "rv32i_m/F/src/flw-align-01.S",
    "rv32i_m/F/src/fmadd_b1-01.S",
    "rv32i_m/F/src/fmadd_b14-01.S",
    "rv32i_m/F/src/fmadd_b15-01.S",
    "rv32i_m/F/src/fmadd_b16-01.S",
    "rv32i_m/F/src/fmadd_b17-01.S",
    "rv32i_m/F/src/fmadd_b18-01.S",
    "rv32i_m/F/src/fmadd_b2-01.S",
    "rv32i_m/F/src/fmadd_b3-01.S",
    "rv32i_m/F/src/fmadd_b4-01.S",
    "rv32i_m/F/src/fmadd_b5-01.S",
    "rv32i_m/F/src/fmadd_b6-01.S",
    "rv32i_m/F/src/fmadd_b7-01.S",
    "rv32i_m/F/src/fmadd_b8-01.S",
    "rv32i_m/F/src/fmax_b1-01.S",
    "rv32i_m/F/src/fmax_b19-01.S",
    "rv32i_m/F/src/fmin_b1-01.S",
    "rv32i_m/F/src/fmin_b19-01.S",
    "rv32i_m/F/src/fmsub_b1-01.S",
    "rv32i_m/F/src/fmsub_b14-01.S",
    //"rv32i_m/F/src/fmsub_b15-01.S",
    "rv32i_m/F/src/fmsub_b16-01.S",
    "rv32i_m/F/src/fmsub_b17-01.S",
    "rv32i_m/F/src/fmsub_b18-01.S",
    "rv32i_m/F/src/fmsub_b2-01.S",
    "rv32i_m/F/src/fmsub_b3-01.S",
    "rv32i_m/F/src/fmsub_b4-01.S",
    "rv32i_m/F/src/fmsub_b5-01.S",
    "rv32i_m/F/src/fmsub_b6-01.S",
    "rv32i_m/F/src/fmsub_b7-01.S",
    "rv32i_m/F/src/fmsub_b8-01.S",
    "rv32i_m/F/src/fmul_b1-01.S",
    "rv32i_m/F/src/fmul_b2-01.S",
    "rv32i_m/F/src/fmul_b3-01.S",
    "rv32i_m/F/src/fmul_b4-01.S",
    "rv32i_m/F/src/fmul_b5-01.S",
    "rv32i_m/F/src/fmul_b6-01.S",
    "rv32i_m/F/src/fmul_b7-01.S",
    "rv32i_m/F/src/fmul_b8-01.S",
    "rv32i_m/F/src/fmul_b9-01.S",
    "rv32i_m/F/src/fmv.w.x_b25-01.S",
    "rv32i_m/F/src/fmv.w.x_b26-01.S",
    "rv32i_m/F/src/fmv.x.w_b1-01.S",
    "rv32i_m/F/src/fmv.x.w_b22-01.S",
    "rv32i_m/F/src/fmv.x.w_b23-01.S",
    "rv32i_m/F/src/fmv.x.w_b24-01.S",
    "rv32i_m/F/src/fmv.x.w_b27-01.S",
    "rv32i_m/F/src/fmv.x.w_b28-01.S",
    "rv32i_m/F/src/fmv.x.w_b29-01.S",
    "rv32i_m/F/src/fnmadd_b1-01.S",
    "rv32i_m/F/src/fnmadd_b14-01.S",
    // "rv32i_m/F/src/fnmadd_b15-01.S",
    "rv32i_m/F/src/fnmadd_b16-01.S",
    "rv32i_m/F/src/fnmadd_b17-01.S",
    "rv32i_m/F/src/fnmadd_b18-01.S",
    "rv32i_m/F/src/fnmadd_b2-01.S",
    "rv32i_m/F/src/fnmadd_b3-01.S",
    "rv32i_m/F/src/fnmadd_b4-01.S",
    "rv32i_m/F/src/fnmadd_b5-01.S",
    "rv32i_m/F/src/fnmadd_b6-01.S",
    "rv32i_m/F/src/fnmadd_b7-01.S",
    "rv32i_m/F/src/fnmadd_b8-01.S",
    "rv32i_m/F/src/fnmsub_b1-01.S",
    "rv32i_m/F/src/fnmsub_b14-01.S",
    // "rv32i_m/F/src/fnmsub_b15-01.S",
    "rv32i_m/F/src/fnmsub_b16-01.S",
    "rv32i_m/F/src/fnmsub_b17-01.S",
    "rv32i_m/F/src/fnmsub_b18-01.S",
    "rv32i_m/F/src/fnmsub_b2-01.S",
    "rv32i_m/F/src/fnmsub_b3-01.S",
    "rv32i_m/F/src/fnmsub_b4-01.S",
    "rv32i_m/F/src/fnmsub_b5-01.S",
    "rv32i_m/F/src/fnmsub_b6-01.S",
    "rv32i_m/F/src/fnmsub_b7-01.S",
    "rv32i_m/F/src/fnmsub_b8-01.S",
    "rv32i_m/F/src/fsgnj_b1-01.S",
    "rv32i_m/F/src/fsgnjn_b1-01.S",
    "rv32i_m/F/src/fsgnjx_b1-01.S",
    "rv32i_m/F/src/fsqrt_b1-01.S",
    "rv32i_m/F/src/fsqrt_b20-01.S",
    "rv32i_m/F/src/fsqrt_b2-01.S",
    "rv32i_m/F/src/fsqrt_b3-01.S",
    "rv32i_m/F/src/fsqrt_b4-01.S",
    "rv32i_m/F/src/fsqrt_b5-01.S",
    "rv32i_m/F/src/fsqrt_b7-01.S",
    "rv32i_m/F/src/fsqrt_b8-01.S",
    "rv32i_m/F/src/fsqrt_b9-01.S",
    "rv32i_m/F/src/fsub_b10-01.S",
    "rv32i_m/F/src/fsub_b1-01.S",
    "rv32i_m/F/src/fsub_b11-01.S",
    "rv32i_m/F/src/fsub_b12-01.S",
    "rv32i_m/F/src/fsub_b13-01.S",
    "rv32i_m/F/src/fsub_b2-01.S",
    "rv32i_m/F/src/fsub_b3-01.S",
    "rv32i_m/F/src/fsub_b4-01.S",
    "rv32i_m/F/src/fsub_b5-01.S",
    "rv32i_m/F/src/fsub_b7-01.S",
    "rv32i_m/F/src/fsub_b8-01.S",
    "rv32i_m/F/src/fsw-align-01.S"
    };

  string arch32d[] = '{
    `RISCVARCHTEST,
    "rv32i_m/D/src/fadd.d_b10-01.S",
    "rv32i_m/D/src/fadd.d_b1-01.S",
    "rv32i_m/D/src/fadd.d_b11-01.S",
    "rv32i_m/D/src/fadd.d_b12-01.S",
    "rv32i_m/D/src/fadd.d_b13-01.S",
    "rv32i_m/D/src/fadd.d_b2-01.S",
    "rv32i_m/D/src/fadd.d_b3-01.S",
    "rv32i_m/D/src/fadd.d_b4-01.S",
    "rv32i_m/D/src/fadd.d_b5-01.S",
    "rv32i_m/D/src/fadd.d_b7-01.S",
    "rv32i_m/D/src/fadd.d_b8-01.S",
    "rv32i_m/D/src/fclass.d_b1-01.S",
    "rv32i_m/D/src/fcvt.d.s_b1-01.S",
    "rv32i_m/D/src/fcvt.d.s_b22-01.S",
    "rv32i_m/D/src/fcvt.d.s_b23-01.S",
    "rv32i_m/D/src/fcvt.d.s_b24-01.S",
    "rv32i_m/D/src/fcvt.d.s_b27-01.S",
    "rv32i_m/D/src/fcvt.d.s_b28-01.S",
    "rv32i_m/D/src/fcvt.d.s_b29-01.S",
    "rv32i_m/D/src/fcvt.d.w_b25-01.S",
    "rv32i_m/D/src/fcvt.d.w_b26-01.S",
    "rv32i_m/D/src/fcvt.d.wu_b25-01.S",
    "rv32i_m/D/src/fcvt.d.wu_b26-01.S",
    "rv32i_m/D/src/fcvt.s.d_b1-01.S",
    "rv32i_m/D/src/fcvt.s.d_b22-01.S",
    "rv32i_m/D/src/fcvt.s.d_b23-01.S",
    "rv32i_m/D/src/fcvt.s.d_b24-01.S",
    "rv32i_m/D/src/fcvt.s.d_b27-01.S",
    "rv32i_m/D/src/fcvt.s.d_b28-01.S",
    "rv32i_m/D/src/fcvt.s.d_b29-01.S",
    "rv32i_m/D/src/fcvt.w.d_b1-01.S",
    "rv32i_m/D/src/fcvt.w.d_b22-01.S",
    "rv32i_m/D/src/fcvt.w.d_b23-01.S",
    "rv32i_m/D/src/fcvt.w.d_b24-01.S",
    "rv32i_m/D/src/fcvt.w.d_b27-01.S",
    "rv32i_m/D/src/fcvt.w.d_b28-01.S",
    "rv32i_m/D/src/fcvt.w.d_b29-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b1-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b22-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b23-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b24-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b27-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b28-01.S",
    "rv32i_m/D/src/fcvt.wu.d_b29-01.S",
    "rv32i_m/D/src/fdiv.d_b1-01.S",
    "rv32i_m/D/src/fdiv.d_b20-01.S",
    "rv32i_m/D/src/fdiv.d_b2-01.S",
    "rv32i_m/D/src/fdiv.d_b21-01.S",
    "rv32i_m/D/src/fdiv.d_b3-01.S",
    "rv32i_m/D/src/fdiv.d_b4-01.S",
    "rv32i_m/D/src/fdiv.d_b5-01.S",
    "rv32i_m/D/src/fdiv.d_b6-01.S",
    "rv32i_m/D/src/fdiv.d_b7-01.S",
    "rv32i_m/D/src/fdiv.d_b8-01.S",
    "rv32i_m/D/src/fdiv.d_b9-01.S",
    "rv32i_m/D/src/feq.d_b1-01.S",
    "rv32i_m/D/src/feq.d_b19-01.S",
    "rv32i_m/D/src/fle.d_b1-01.S",
    "rv32i_m/D/src/fle.d_b19-01.S",
    "rv32i_m/D/src/flt.d_b1-01.S",
    "rv32i_m/D/src/flt.d_b19-01.S",
    "rv32i_m/D/src/fld-align-01.S", 
    "rv32i_m/D/src/fsd-align-01.S", 
    "rv32i_m/D/src/fmadd.d_b14-01.S",
    "rv32i_m/D/src/fmadd.d_b16-01.S",
    "rv32i_m/D/src/fmadd.d_b17-01.S",
    "rv32i_m/D/src/fmadd.d_b18-01.S",
    "rv32i_m/D/src/fmadd.d_b2-01.S",
    "rv32i_m/D/src/fmadd.d_b3-01.S",
    "rv32i_m/D/src/fmadd.d_b4-01.S",
    "rv32i_m/D/src/fmadd.d_b5-01.S",
    "rv32i_m/D/src/fmadd.d_b6-01.S",
    "rv32i_m/D/src/fmadd.d_b7-01.S",
    "rv32i_m/D/src/fmadd.d_b8-01.S",
    "rv32i_m/D/src/fmax.d_b1-01.S",
    "rv32i_m/D/src/fmax.d_b19-01.S",
    "rv32i_m/D/src/fmin.d_b1-01.S",
    "rv32i_m/D/src/fmin.d_b19-01.S",
    "rv32i_m/D/src/fmsub.d_b14-01.S",
    "rv32i_m/D/src/fmsub.d_b16-01.S",
    "rv32i_m/D/src/fmsub.d_b17-01.S",
    "rv32i_m/D/src/fmsub.d_b18-01.S",
    "rv32i_m/D/src/fmsub.d_b2-01.S",
    "rv32i_m/D/src/fmsub.d_b3-01.S",
    "rv32i_m/D/src/fmsub.d_b4-01.S",
    "rv32i_m/D/src/fmsub.d_b5-01.S",
    "rv32i_m/D/src/fmsub.d_b6-01.S",
    "rv32i_m/D/src/fmsub.d_b7-01.S",
    "rv32i_m/D/src/fmsub.d_b8-01.S",
    "rv32i_m/D/src/fmul.d_b1-01.S",
    "rv32i_m/D/src/fmul.d_b2-01.S",
    "rv32i_m/D/src/fmul.d_b3-01.S",
    "rv32i_m/D/src/fmul.d_b4-01.S",
    "rv32i_m/D/src/fmul.d_b5-01.S",
    "rv32i_m/D/src/fmul.d_b6-01.S",
    "rv32i_m/D/src/fmul.d_b7-01.S",
    "rv32i_m/D/src/fmul.d_b8-01.S",
    "rv32i_m/D/src/fmul.d_b9-01.S",
    "rv32i_m/D/src/fnmadd.d_b14-01.S",
    "rv32i_m/D/src/fnmadd.d_b16-01.S",
    "rv32i_m/D/src/fnmadd.d_b17-01.S",
    "rv32i_m/D/src/fnmadd.d_b18-01.S",
    "rv32i_m/D/src/fnmadd.d_b2-01.S",
    "rv32i_m/D/src/fnmadd.d_b3-01.S",
    "rv32i_m/D/src/fnmadd.d_b4-01.S",
    "rv32i_m/D/src/fnmadd.d_b5-01.S",
    "rv32i_m/D/src/fnmadd.d_b6-01.S",
    "rv32i_m/D/src/fnmadd.d_b7-01.S",
    "rv32i_m/D/src/fnmadd.d_b8-01.S",
    "rv32i_m/D/src/fnmsub.d_b14-01.S",
    "rv32i_m/D/src/fnmsub.d_b16-01.S",
    "rv32i_m/D/src/fnmsub.d_b17-01.S",
    "rv32i_m/D/src/fnmsub.d_b18-01.S",
    "rv32i_m/D/src/fnmsub.d_b2-01.S",
    "rv32i_m/D/src/fnmsub.d_b3-01.S",
    "rv32i_m/D/src/fnmsub.d_b4-01.S",
    "rv32i_m/D/src/fnmsub.d_b5-01.S",
    "rv32i_m/D/src/fnmsub.d_b6-01.S",
    "rv32i_m/D/src/fnmsub.d_b7-01.S",
    "rv32i_m/D/src/fnmsub.d_b8-01.S",
    "rv32i_m/D/src/fsgnj.d_b1-01.S",
    "rv32i_m/D/src/fsgnjn.d_b1-01.S",
    "rv32i_m/D/src/fsgnjx.d_b1-01.S",
    "rv32i_m/D/src/fsqrt.d_b1-01.S",
    "rv32i_m/D/src/fsqrt.d_b20-01.S",
    "rv32i_m/D/src/fsqrt.d_b2-01.S",
    "rv32i_m/D/src/fsqrt.d_b3-01.S",
    "rv32i_m/D/src/fsqrt.d_b4-01.S",
    "rv32i_m/D/src/fsqrt.d_b5-01.S",
    "rv32i_m/D/src/fsqrt.d_b7-01.S",
    "rv32i_m/D/src/fsqrt.d_b8-01.S",
    "rv32i_m/D/src/fsqrt.d_b9-01.S",
    "rv32i_m/D/src/fssub.d_b10-01.S",
    "rv32i_m/D/src/fssub.d_b1-01.S",
    "rv32i_m/D/src/fssub.d_b11-01.S",
    "rv32i_m/D/src/fssub.d_b12-01.S",
    "rv32i_m/D/src/fssub.d_b13-01.S",
    "rv32i_m/D/src/fssub.d_b2-01.S",
    "rv32i_m/D/src/fssub.d_b3-01.S",
    "rv32i_m/D/src/fssub.d_b4-01.S",
    "rv32i_m/D/src/fssub.d_b5-01.S",
    "rv32i_m/D/src/fssub.d_b7-01.S",
    "rv32i_m/D/src/fssub.d_b8-01.S"
};


  string arch32c[] = '{
    `RISCVARCHTEST,
    "rv32i_m/C/src/cadd-01.S",
  "rv32i_m/C/src/caddi-01.S",
  "rv32i_m/C/src/caddi16sp-01.S",
  "rv32i_m/C/src/caddi4spn-01.S",
  "rv32i_m/C/src/cand-01.S",
  "rv32i_m/C/src/candi-01.S",
  "rv32i_m/C/src/cbeqz-01.S",
  "rv32i_m/C/src/cbnez-01.S",
  "rv32i_m/C/src/cj-01.S",
  "rv32i_m/C/src/cjal-01.S",
  "rv32i_m/C/src/cjalr-01.S",
  "rv32i_m/C/src/cjr-01.S",
  "rv32i_m/C/src/cli-01.S",
  "rv32i_m/C/src/clui-01.S",
  "rv32i_m/C/src/clw-01.S",
  "rv32i_m/C/src/clwsp-01.S",
  "rv32i_m/C/src/cmv-01.S",
  "rv32i_m/C/src/cnop-01.S",
  "rv32i_m/C/src/cor-01.S",
  "rv32i_m/C/src/cslli-01.S",
  "rv32i_m/C/src/csrai-01.S",
  "rv32i_m/C/src/csrli-01.S",
  "rv32i_m/C/src/csub-01.S",
  "rv32i_m/C/src/csw-01.S",
  "rv32i_m/C/src/cswsp-01.S",
  "rv32i_m/C/src/cxor-01.S"
  };

  string arch32cpriv[] = '{
  //  `RISCVARCHTEST,
  "rv32i_m/C/src/cebreak-01.S"
  };      


  string arch32i[] = '{
    `RISCVARCHTEST,
    "rv32i_m/I/src/add-01.S",
    "rv32i_m/I/src/addi-01.S",
    "rv32i_m/I/src/and-01.S",
    "rv32i_m/I/src/andi-01.S",
    "rv32i_m/I/src/auipc-01.S",
    "rv32i_m/I/src/beq-01.S",
    "rv32i_m/I/src/bge-01.S",
    "rv32i_m/I/src/bgeu-01.S",
    "rv32i_m/I/src/blt-01.S",
    "rv32i_m/I/src/bltu-01.S",
    "rv32i_m/I/src/bne-01.S",
    "rv32i_m/I/src/fence-01.S",
    "rv32i_m/I/src/jal-01.S",
    "rv32i_m/I/src/jalr-01.S",
    "rv32i_m/I/src/lb-align-01.S",
    "rv32i_m/I/src/lbu-align-01.S",
    "rv32i_m/I/src/lh-align-01.S",
    "rv32i_m/I/src/lhu-align-01.S",
    "rv32i_m/I/src/lui-01.S",
    "rv32i_m/I/src/lw-align-01.S",
    "rv32i_m/I/src/or-01.S",
    "rv32i_m/I/src/ori-01.S",
    "rv32i_m/I/src/sb-align-01.S",
    "rv32i_m/I/src/sh-align-01.S",
    "rv32i_m/I/src/sll-01.S",
    "rv32i_m/I/src/slli-01.S",
    "rv32i_m/I/src/slt-01.S",
    "rv32i_m/I/src/slti-01.S",
    "rv32i_m/I/src/sltiu-01.S",
    "rv32i_m/I/src/sltu-01.S",
    "rv32i_m/I/src/sra-01.S",
    "rv32i_m/I/src/srai-01.S",
    "rv32i_m/I/src/srl-01.S",
    "rv32i_m/I/src/srli-01.S",
    "rv32i_m/I/src/sub-01.S",
    "rv32i_m/I/src/sw-align-01.S",
    "rv32i_m/I/src/xor-01.S",
    "rv32i_m/I/src/xori-01.S"
  };

 string wally64i[] = '{
    `WALLYTEST,
    "rv64i_m/I/src/WALLY-ADD.S",
    "rv64i_m/I/src/WALLY-SLT.S",
    "rv64i_m/I/src/WALLY-SLTU.S",
    "rv64i_m/I/src/WALLY-SUB.S",
    "rv64i_m/I/src/WALLY-XOR.S"
 };

 
 string wally64priv[] = '{
    `WALLYTEST,
//    "rv64i_m/privilege/src/BUG66",
    "rv64i_m/privilege/src/WALLY-csr-permission-s-01.S",
    "rv64i_m/privilege/src/WALLY-csr-permission-u-01.S",
    "rv64i_m/privilege/src/WALLY-mie-01.S",
    "rv64i_m/privilege/src/WALLY-minfo-01.S",
    "rv64i_m/privilege/src/WALLY-misa-01.S",
    "rv64i_m/privilege/src/WALLY-mmu-sv39-01.S",
    "rv64i_m/privilege/src/WALLY-mmu-sv48-01.S",
    "rv64i_m/privilege/src/WALLY-mtvec-01.S",
    "rv64i_m/privilege/src/WALLY-pma-01.S",
    "rv64i_m/privilege/src/WALLY-pmp-01.S",
    "rv64i_m/privilege/src/WALLY-sie-01.S",
    "rv64i_m/privilege/src/WALLY-status-mie-01.S",
    "rv64i_m/privilege/src/WALLY-status-sie-01.S",
    "rv64i_m/privilege/src/WALLY-status-tw-01.S",
    "rv64i_m/privilege/src/WALLY-status-tvm-01.S",
    "rv64i_m/privilege/src/WALLY-status-fp-enabled-01.S",
    "rv64i_m/privilege/src/WALLY-stvec-01.S",
    "rv64i_m/privilege/src/WALLY-trap-01.S",
    "rv64i_m/privilege/src/WALLY-trap-s-01.S",
    "rv64i_m/privilege/src/WALLY-trap-sret-01.S",
    "rv64i_m/privilege/src/WALLY-trap-u-01.S",
    "rv64i_m/privilege/src/WALLY-wfi-01.S",
    "rv64i_m/privilege/src/WALLY-endianness-01.S",
    "rv64i_m/privilege/src/WALLY-status-xlen-01.S",
    "rv64i_m/privilege/src/WALLY-satp-invalid-01.S"
 };

 string wally64periph[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/src/WALLY-periph-01.S",
    "rv64i_m/privilege/src/WALLY-clint-01.S",
    "rv64i_m/privilege/src/WALLY-gpio-01.S",
    "rv64i_m/privilege/src/WALLY-plic-01.S",
    "rv64i_m/privilege/src/WALLY-plic-s-01.S",
    "rv64i_m/privilege/src/WALLY-uart-01.S"
 };

 string wally32e[] = '{
    `WALLYTEST,
    "rv32i_m/I/src/E-add-01.S",
    "rv32i_m/I/src/E-addi-01.S",
    "rv32i_m/I/src/E-and-01.S",
    "rv32i_m/I/src/E-andi-01.S",
    "rv32i_m/I/src/E-auipc-01.S",
    "rv32i_m/I/src/E-bge-01.S",
    "rv32i_m/I/src/E-bgeu-01.S",
    "rv32i_m/I/src/E-blt-01.S",
    "rv32i_m/I/src/E-bltu-01.S",
    "rv32i_m/I/src/E-bne-01.S",
    "rv32i_m/I/src/E-jal-01.S",
    "rv32i_m/I/src/E-jalr-01.S",
    "rv32i_m/I/src/E-lb-align-01.S",
    "rv32i_m/I/src/E-lbu-align-01.S",
    "rv32i_m/I/src/E-lh-align-01.S",
    "rv32i_m/I/src/E-lhu-align-01.S",
    "rv32i_m/I/src/E-lui-01.S",
    "rv32i_m/I/src/E-lw-align-01.S",
    "rv32i_m/I/src/E-or-01.S",
    "rv32i_m/I/src/E-ori-01.S",
    "rv32i_m/I/src/E-sb-align-01.S",
    "rv32i_m/I/src/E-sh-align-01.S",
    "rv32i_m/I/src/E-sll-01.S",
    "rv32i_m/I/src/E-slli-01.S",
    "rv32i_m/I/src/E-slt-01.S",
    "rv32i_m/I/src/E-slti-01.S",
    "rv32i_m/I/src/E-sltiu-01.S",
    "rv32i_m/I/src/E-sltu-01.S",
    "rv32i_m/I/src/E-sra-01.S",
    "rv32i_m/I/src/E-srai-01.S",
    "rv32i_m/I/src/E-srl-01.S",
    "rv32i_m/I/src/E-srli-01.S",
    "rv32i_m/I/src/E-sub-01.S",
    "rv32i_m/I/src/E-sw-align-01.S",
    "rv32i_m/I/src/E-xor-01.S",
    "rv32i_m/I/src/E-xori-01.S"
 };

 string wally32i[] = '{
    `WALLYTEST,
    "rv32i_m/I/src/WALLY-ADD.S",
    "rv32i_m/I/src/WALLY-SLT.S",
    "rv32i_m/I/src/WALLY-SLTU.S",
    "rv32i_m/I/src/WALLY-SUB.S",
    "rv32i_m/I/src/WALLY-XOR.S" 
 };


 string wally32priv[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/src/WALLY-csr-permission-s-01.S",
    "rv32i_m/privilege/src/WALLY-csr-permission-u-01.S",
    "rv32i_m/privilege/src/WALLY-mie-01.S",
    "rv32i_m/privilege/src/WALLY-minfo-01.S",
    "rv32i_m/privilege/src/WALLY-misa-01.S",
    "rv32i_m/privilege/src/WALLY-mmu-sv32-01.S",
    "rv32i_m/privilege/src/WALLY-mtvec-01.S",
    "rv32i_m/privilege/src/WALLY-pma-01.S",
    "rv32i_m/privilege/src/WALLY-pmp-01.S",
    "rv32i_m/privilege/src/WALLY-sie-01.S",
    "rv32i_m/privilege/src/WALLY-status-mie-01.S",
    "rv32i_m/privilege/src/WALLY-status-sie-01.S",
    "rv32i_m/privilege/src/WALLY-status-tw-01.S",
    "rv32i_m/privilege/src/WALLY-status-tvm-01.S",
    "rv32i_m/privilege/src/WALLY-status-fp-enabled-01.S",
    "rv32i_m/privilege/src/WALLY-stvec-01.S",
    "rv32i_m/privilege/src/WALLY-trap-01.S",
    "rv32i_m/privilege/src/WALLY-trap-s-01.S",
    "rv32i_m/privilege/src/WALLY-trap-sret-01.S",
    "rv32i_m/privilege/src/WALLY-trap-u-01.S",
    "rv32i_m/privilege/src/WALLY-wfi-01.S",
    "rv32i_m/privilege/src/WALLY-endianness-01.S",
    "rv32i_m/privilege/src/WALLY-satp-invalid-01.S"
 };

 string wally32periph[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/src/WALLY-periph-01.S",
    "rv32i_m/privilege/src/WALLY-gpio-01.S",
    "rv32i_m/privilege/src/WALLY-clint-01.S",
    "rv32i_m/privilege/src/WALLY-uart-01.S",
    "rv32i_m/privilege/src/WALLY-plic-01.S",
    "rv32i_m/privilege/src/WALLY-plic-s-01.S"
 };


 string wally32d[] = '{
    `WALLYTEST,
    "rv32i_m/D/src/WALLY-fld-01.S"
 };

 string fpga[] = '{
    `CUSTOM,
    "NULL"
 };

 string custom[] = '{
    `CUSTOM,
    "debug",
    "simple",
    "cacheTest"
 };
  string testsBP64[] = '{
    `IMPERASTEST,
    "rv64BP/simple"
//    "rv64BP/mmm",
//    "rv64BP/linpack_bench",
//    "rv64BP/sieve",
//    "rv64BP/qsort",
//    "rv64BP/dhrystone"
  };


 string ahb[] = '{
    `RISCVARCHTEST,
    "rv64i_m/F/src/fadd_b11-01.S"
 };

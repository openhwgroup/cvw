///////////////////////////////////////////
// bsg_dmc_config_apb.sv
//
// Written: infinitymdm@gmail.com 3 June 2024
//
// Purpose: Synchronized configuration registers for BSG memory controller
// 
// Documentation: 
//
// A component of the CORE-V-WALLY configurable RISC-V project.
// https://github.com/openhwgroup/cvw
// 
// Copyright (C) 2021-24 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

module bsg_dmc_config_apb #(parameter APB_DATA_SIZE = 64) (
  input  logic                     PCLK, PRESETn,
  input  logic                     PSEL,
  input  logic [7:0]               PADDR,
  input  logic [APB_DATA_SIZE-1:0] PWDATA,
  input  logic                     PWRITE,
  input  logic                     PENABLE,
  output logic [APB_DATA_SIZE-1:0] PRDATA,
  output logic                     PREADY,
  input  logic                     ui_clk,
  output logic [15:0]              dmc_trefi,
  output logic [3:0]               dmc_tmrd,
  output logic [3:0]               dmc_trfc,
  output logic [3:0]               dmc_trc,
  output logic [3:0]               dmc_trp,
  output logic [3:0]               dmc_tras,
  output logic [3:0]               dmc_trrd,
  output logic [3:0]               dmc_trcd,
  output logic [3:0]               dmc_twr,
  output logic [3:0]               dmc_twtr,
  output logic [3:0]               dmc_trtp,
  output logic [3:0]               dmc_tcas,
  output logic [3:0]               dmc_col_width,
  output logic [3:0]               dmc_row_width,
  output logic [1:0]               dmc_bank_width,
  output logic [5:0]               dmc_bank_pos,
  output logic [2:0]               dmc_dqs_sel_cal,
  output logic [15:0]              dmc_init_cycles,
  output logic                     dmc_config_changed
);

  logic [7:0]   entry, wentry;
  logic         wren;
  logic [15:0]  wdata;
  logic [15:0]  rdata;
  logic         fifo_full, fifo_deq;

  assign entry  = {PADDR[7:3], 3'b0};
  assign PREADY = ~fifo_full;

  // Send writes to ui_clk domain
  assign wren = PWRITE & PENABLE & PSEL;
  bsg_async_fifo #(
    .lg_size_p(3),
    .width_p(8 + 16) // entry + data
  ) dmc_config_fifo (
    .w_clk_i(PCLK),
    .w_reset_i(~PRESETn),
    .w_enq_i(wren),
    .w_data_i({entry, PWDATA[15:0]}),
    .w_full_o(fifo_full),
    .r_clk_i(ui_clk),
    .r_reset_i(~PRESETn),
    .r_deq_i(fifo_deq & dmc_config_changed),
    .r_data_o({wentry, wdata}),
    .r_valid_o(dmc_config_changed)
  );
  flopr #(1) deqreg (ui_clk, ~PRESETn, dmc_config_changed, fifo_deq);

  // Write on ui_clk with async reset
  always_ff @(posedge ui_clk, negedge PRESETn) begin
    if (~PRESETn) begin
      // TODO: Should these be reset to Micron defaults instead?
      dmc_trefi        <= 0;
      dmc_tmrd         <= 0;
      dmc_trfc         <= 0;
      dmc_trc          <= 0;
      dmc_trp          <= 0;
      dmc_tras         <= 0;
      dmc_trrd         <= 0;
      dmc_trcd         <= 0;
      dmc_twr          <= 0;
      dmc_twtr         <= 0;
      dmc_trtp         <= 0;
      dmc_tcas         <= 0;
      dmc_col_width    <= 0;
      dmc_row_width    <= 0;
      dmc_bank_width   <= 0;
      dmc_bank_pos     <= 0;
      dmc_dqs_sel_cal  <= 0;
      dmc_init_cycles  <= 0;
    end else begin
      if (dmc_config_changed) begin
        case (wentry)
          8'h00: dmc_trefi       <= wdata;
          8'h08: dmc_tmrd        <= wdata[3:0];
          8'h10: dmc_trfc        <= wdata[3:0];
          8'h18: dmc_trc         <= wdata[3:0];
          8'h20: dmc_trp         <= wdata[3:0];
          8'h28: dmc_tras        <= wdata[3:0];
          8'h30: dmc_trrd        <= wdata[3:0];
          8'h38: dmc_trcd        <= wdata[3:0];
          8'h40: dmc_twr         <= wdata[3:0];
          8'h48: dmc_twtr        <= wdata[3:0];
          8'h50: dmc_trtp        <= wdata[3:0];
          8'h58: dmc_tcas        <= wdata[3:0];
          8'h60: dmc_col_width   <= wdata[3:0];
          8'h68: dmc_row_width   <= wdata[3:0];
          8'h70: dmc_bank_width  <= wdata[1:0];
          8'h78: dmc_bank_pos    <= wdata[5:0];
          8'h80: dmc_dqs_sel_cal <= wdata[2:0];
          8'h88: dmc_init_cycles <= wdata;
        endcase
      end
    end
  end

  // Read on PCLK
  assign PRDATA = {{APB_DATA_SIZE-17{1'b0}}, rdata};
  always_ff @(posedge PCLK) begin
    case (entry)
      8'h00:   rdata <=         dmc_trefi;
      8'h08:   rdata <= {12'b0, dmc_tmrd};
      8'h10:   rdata <= {12'b0, dmc_trfc};
      8'h18:   rdata <= {12'b0, dmc_trc};
      8'h20:   rdata <= {12'b0, dmc_trp};
      8'h28:   rdata <= {12'b0, dmc_tras};
      8'h30:   rdata <= {12'b0, dmc_trrd};
      8'h38:   rdata <= {12'b0, dmc_trcd};
      8'h40:   rdata <= {12'b0, dmc_twr};
      8'h48:   rdata <= {12'b0, dmc_twtr};
      8'h50:   rdata <= {12'b0, dmc_trtp};
      8'h58:   rdata <= {12'b0, dmc_tcas};
      8'h60:   rdata <= {12'b0, dmc_col_width};
      8'h68:   rdata <= {12'b0, dmc_row_width};
      8'h70:   rdata <= {14'b0, dmc_bank_width};
      8'h78:   rdata <= {10'b0, dmc_bank_pos};
      8'h80:   rdata <= {13'b0, dmc_dqs_sel_cal};
      8'h88:   rdata <=         dmc_init_cycles;
      default: rdata <= 0;
    endcase
  end

endmodule

///////////////////////////////////////////
// tests.vh
//
// Written: David_Harris@hmc.edu 7 October 2021
// Modified: 
//
// Purpose: List of tests to apply
// 
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, 
// modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software 
// is furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES 
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS 
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT 
// OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
///////////////////////////////////////////

`define IMPERASTEST   "0"
`define RISCVARCHTEST "1"
`define WALLYTEST "2"
`define MYIMPERASTEST   "3"
`define COREMARK "4"
// *** remove MYIMPERASTEST cases when ported 

string tvpaths[] = '{
    "../../addins/imperas-riscv-tests/work/",
    "../../addins/riscv-arch-test/work/",
    "../../tests/wally-riscv-arch-test/work/",
    "../../tests/imperas-riscv-tests/work/",
    "../../benchmarks/riscv-coremark/work/"
};

   // *** make sure these are somewhere
  string coremark[] = '{
    `COREMARK,
    "coremark.bare.riscv", "100000"
  };

  string wally64a[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-AMO", "2210",
    "rv64i_m/privilege/WALLY-LRSC", "2410"
  };

    string wally32a[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/WALLY-AMO", "2310",
    "rv32i_m/privilege/WALLY-LRSC", "2310"
  };

  // *** restore CSR tests from Imperas old

    string extra64i[] = '{
    `MYIMPERASTEST,
    "rv64i_m/I/WALLY-ADD", "4000",
    "rv64i_m/I/WALLY-SUB", "4000",
    "rv64i_m/I/WALLY-ADDI", "3000",
    "rv64i_m/I/WALLY-ANDI", "3000",
    "rv64i_m/I/WALLY-ORI", "3000",
    "rv64i_m/I/WALLY-XORI", "3000",
    "rv64i_m/I/WALLY-SLTI", "3000",
    "rv64i_m/I/WALLY-SLTIU", "3000",
    "rv64i_m/I/WALLY-SLLI", "3000",
    "rv64i_m/I/WALLY-SRLI", "3000",
    "rv64i_m/I/WALLY-SRAI", "3000",
    "rv64i_m/I/WALLY-JAL", "4000",
    "rv64i_m/I/WALLY-JALR", "3000",
    "rv64i_m/I/WALLY-STORE", "3000",
    "rv64i_m/I/WALLY-ADDIW", "3000",
    "rv64i_m/I/WALLY-SLLIW", "3000",
    "rv64i_m/I/WALLY-SRLIW", "3000",
    "rv64i_m/I/WALLY-SRAIW", "3000",
    "rv64i_m/I/WALLY-ADDW", "4000",
    "rv64i_m/I/WALLY-SUBW", "4000",
    "rv64i_m/I/WALLY-SLLW", "3000",
    "rv64i_m/I/WALLY-SRLW", "3000",
    "rv64i_m/I/WALLY-SRAW", "3000",
    "rv64i_m/I/WALLY-BEQ" ,"5000",
    "rv64i_m/I/WALLY-BNE", "5000 ",
    "rv64i_m/I/WALLY-BLTU", "5000 ",
    "rv64i_m/I/WALLY-BLT", "5000",
    "rv64i_m/I/WALLY-BGE", "5000 ",
    "rv64i_m/I/WALLY-BGEU", "5000 ",
    "rv64i_m/I/WALLY-CSRRW", "4000",
    "rv64i_m/I/WALLY-CSRRS", "4000",
    "rv64i_m/I/WALLY-CSRRC", "5000",
    "rv64i_m/I/WALLY-CSRRWI", "4000",
    "rv64i_m/I/WALLY-CSRRSI", "4000",
    "rv64i_m/I/WALLY-CSRRCI", "4000" 
  };

  
string imperas32f[] = '{
    `IMPERASTEST,
    "rv32i_m/F/FADD-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FADD-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FADD-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FADD-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FADD-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FADD-S-RDN-01", "002010",
    "rv32i_m/F/FADD-S-RMM-01", "002010",
    "rv32i_m/F/FADD-S-RNE-01", "002010",
    "rv32i_m/F/FADD-S-RTZ-01", "002010",
    "rv32i_m/F/FADD-S-RUP-01", "002010",
    "rv32i_m/F/FCLASS-S-01", "002010",
    "rv32i_m/F/FCVT-S-W-DYN-RDN-01", "002010",
    "rv32i_m/F/FCVT-S-W-DYN-RMM-01", "002010",
    "rv32i_m/F/FCVT-S-W-DYN-RNE-01", "002010",
    "rv32i_m/F/FCVT-S-W-DYN-RTZ-01", "002010",
    "rv32i_m/F/FCVT-S-W-DYN-RUP-01", "002010",
    "rv32i_m/F/FCVT-S-W-RDN-01", "002010",
    "rv32i_m/F/FCVT-S-W-RMM-01", "002010",
    "rv32i_m/F/FCVT-S-W-RNE-01", "002010",
    "rv32i_m/F/FCVT-S-W-RTZ-01", "002010",
    "rv32i_m/F/FCVT-S-W-RUP-01", "002010",
    "rv32i_m/F/FCVT-S-WU-DYN-RDN-01", "002010",
    "rv32i_m/F/FCVT-S-WU-DYN-RMM-01", "002010",
    "rv32i_m/F/FCVT-S-WU-DYN-RNE-01", "002010",
    "rv32i_m/F/FCVT-S-WU-DYN-RTZ-01", "002010",
    "rv32i_m/F/FCVT-S-WU-DYN-RUP-01", "002010",
    "rv32i_m/F/FCVT-S-WU-RDN-01", "002010",
    "rv32i_m/F/FCVT-S-WU-RMM-01", "002010",
    "rv32i_m/F/FCVT-S-WU-RNE-01", "002010",
    "rv32i_m/F/FCVT-S-WU-RTZ-01", "002010",
    "rv32i_m/F/FCVT-S-WU-RUP-01", "002010",
    "rv32i_m/F/FCVT-W-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FCVT-W-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FCVT-W-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FCVT-W-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FCVT-W-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FCVT-W-S-RDN-01", "002010",
    "rv32i_m/F/FCVT-W-S-RMM-01", "002010",
    "rv32i_m/F/FCVT-W-S-RNE-01", "002010",
    "rv32i_m/F/FCVT-W-S-RTZ-01", "002010",
    "rv32i_m/F/FCVT-W-S-RUP-01", "002010",
    "rv32i_m/F/FCVT-WU-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FCVT-WU-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FCVT-WU-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FCVT-WU-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FCVT-WU-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FCVT-WU-S-RDN-01", "002010",
    "rv32i_m/F/FCVT-WU-S-RMM-01", "002010",
    "rv32i_m/F/FCVT-WU-S-RNE-01", "002010",
    "rv32i_m/F/FCVT-WU-S-RTZ-01", "002010",
    "rv32i_m/F/FCVT-WU-S-RUP-01", "002010",
    // "rv32i_m/F/FDIV-S-DYN-RDN-01", "002010",
    // "rv32i_m/F/FDIV-S-DYN-RMM-01", "002010",
    // "rv32i_m/F/FDIV-S-DYN-RNE-01", "002010",
    // "rv32i_m/F/FDIV-S-DYN-RTZ-01", "002010",
    // "rv32i_m/F/FDIV-S-DYN-RUP-01", "002010",
    // "rv32i_m/F/FDIV-S-RDN-01", "002010",
    // "rv32i_m/F/FDIV-S-RMM-01", "002010",
    // "rv32i_m/F/FDIV-S-RNE-01", "002010",
    // "rv32i_m/F/FDIV-S-RTZ-01", "002010",
    // "rv32i_m/F/FDIV-S-RUP-01", "002010",
    "rv32i_m/F/FEQ-S-01", "002010",
    "rv32i_m/F/FLE-S-01", "002010",
    "rv32i_m/F/FLT-S-01", "002010",
    "rv32i_m/F/FLW-01", "002120",
    "rv32i_m/F/FMADD-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FMADD-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FMADD-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FMADD-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FMADD-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FMADD-S-RDN-01", "002010",
    "rv32i_m/F/FMADD-S-RMM-01", "002010",
    "rv32i_m/F/FMADD-S-RNE-01", "002010",
    "rv32i_m/F/FMADD-S-RTZ-01", "002010",
    "rv32i_m/F/FMADD-S-RUP-01", "002010",
    "rv32i_m/F/FMAX-S-01", "002010",
    "rv32i_m/F/FMIN-S-01", "002010",
    "rv32i_m/F/FMSUB-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FMSUB-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FMSUB-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FMSUB-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FMSUB-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FMSUB-S-RDN-01", "002010",
    "rv32i_m/F/FMSUB-S-RMM-01", "002010",
    "rv32i_m/F/FMSUB-S-RNE-01", "002010",
    "rv32i_m/F/FMSUB-S-RTZ-01", "002010",
    "rv32i_m/F/FMSUB-S-RUP-01", "002010",
    "rv32i_m/F/FMUL-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FMUL-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FMUL-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FMUL-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FMUL-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FMUL-S-RDN-01", "002010",
    "rv32i_m/F/FMUL-S-RMM-01", "002010",
    "rv32i_m/F/FMUL-S-RNE-01", "002010",
    "rv32i_m/F/FMUL-S-RTZ-01", "002010",
    "rv32i_m/F/FMUL-S-RUP-01", "002010",
    "rv32i_m/F/FMV-W-X-01", "002010",
    "rv32i_m/F/FMV-X-W-01", "002010",
    "rv32i_m/F/FNMADD-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FNMADD-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FNMADD-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FNMADD-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FNMADD-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FNMADD-S-RDN-01", "002010",
    "rv32i_m/F/FNMADD-S-RMM-01", "002010",
    "rv32i_m/F/FNMADD-S-RNE-01", "002010",
    "rv32i_m/F/FNMADD-S-RTZ-01", "002010",
    "rv32i_m/F/FNMADD-S-RUP-01", "002010",
    "rv32i_m/F/FNMSUB-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FNMSUB-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FNMSUB-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FNMSUB-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FNMSUB-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FNMSUB-S-RDN-01", "002010",
    "rv32i_m/F/FNMSUB-S-RMM-01", "002010",
    "rv32i_m/F/FNMSUB-S-RNE-01", "002010",
    "rv32i_m/F/FNMSUB-S-RTZ-01", "002010",
    "rv32i_m/F/FNMSUB-S-RUP-01", "002010",
    "rv32i_m/F/FSGNJN-S-01", "002010",
    "rv32i_m/F/FSGNJ-S-01", "002010",
    "rv32i_m/F/FSGNJX-S-01", "002010",
    // "rv32i_m/F/FSQRT-S-DYN-RDN-01", "002010",
    // "rv32i_m/F/FSQRT-S-DYN-RMM-01", "002010",
    // "rv32i_m/F/FSQRT-S-DYN-RNE-01", "002010",
    // "rv32i_m/F/FSQRT-S-DYN-RTZ-01", "002010",
    // "rv32i_m/F/FSQRT-S-DYN-RUP-01", "002010",
    // "rv32i_m/F/FSQRT-S-RDN-01", "002010",
    // "rv32i_m/F/FSQRT-S-RMM-01", "002010",
    // "rv32i_m/F/FSQRT-S-RNE-01", "002010",
    // "rv32i_m/F/FSQRT-S-RTZ-01", "002010",
    // "rv32i_m/F/FSQRT-S-RUP-01", "002010",
    "rv32i_m/F/FSUB-S-DYN-RDN-01", "002010",
    "rv32i_m/F/FSUB-S-DYN-RMM-01", "002010",
    "rv32i_m/F/FSUB-S-DYN-RNE-01", "002010",
    "rv32i_m/F/FSUB-S-DYN-RTZ-01", "002010",
    "rv32i_m/F/FSUB-S-DYN-RUP-01", "002010",
    "rv32i_m/F/FSUB-S-RDN-01", "002010",
    "rv32i_m/F/FSUB-S-RMM-01", "002010",
    "rv32i_m/F/FSUB-S-RNE-01", "002010",
    "rv32i_m/F/FSUB-S-RTZ-01", "002010",
    "rv32i_m/F/FSUB-S-RUP-01", "002010",
    "rv32i_m/F/FSW-01", "002010"
  };

  string imperas64f[] = '{
    `IMPERASTEST,
    "rv64i_m/F/FADD-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FADD-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FADD-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FADD-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FADD-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FADD-S-RDN-01", "002010",
    "rv64i_m/F/FADD-S-RMM-01", "002010",
    "rv64i_m/F/FADD-S-RNE-01", "002010",
    "rv64i_m/F/FADD-S-RTZ-01", "002010",
    "rv64i_m/F/FADD-S-RUP-01", "002010",
    "rv64i_m/F/FCLASS-S-01", "002010",
    "rv64i_m/F/FCVT-L-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-L-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-L-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-L-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-L-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-L-S-RDN-01", "002010",
    "rv64i_m/F/FCVT-L-S-RMM-01", "002010",
    "rv64i_m/F/FCVT-L-S-RNE-01", "002010",
    "rv64i_m/F/FCVT-L-S-RTZ-01", "002010",
    "rv64i_m/F/FCVT-L-S-RUP-01", "002010",
    "rv64i_m/F/FCVT-LU-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-LU-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-LU-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-LU-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-LU-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-LU-S-RDN-01", "002010",
    "rv64i_m/F/FCVT-LU-S-RMM-01", "002010",
    "rv64i_m/F/FCVT-LU-S-RNE-01", "002010",
    "rv64i_m/F/FCVT-LU-S-RTZ-01", "002010",
    "rv64i_m/F/FCVT-LU-S-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-L-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-L-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-L-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-L-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-L-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-L-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-L-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-L-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-L-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-L-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-LU-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-LU-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-LU-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-LU-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-LU-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-LU-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-LU-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-LU-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-LU-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-LU-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-W-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-W-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-W-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-W-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-W-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-W-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-W-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-W-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-W-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-W-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-WU-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-WU-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-WU-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-WU-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-WU-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-S-WU-RDN-01", "002010",
    "rv64i_m/F/FCVT-S-WU-RMM-01", "002010",
    "rv64i_m/F/FCVT-S-WU-RNE-01", "002010",
    "rv64i_m/F/FCVT-S-WU-RTZ-01", "002010",
    "rv64i_m/F/FCVT-S-WU-RUP-01", "002010",
    "rv64i_m/F/FCVT-W-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-W-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-W-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-W-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-W-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-W-S-RDN-01", "002010",
    "rv64i_m/F/FCVT-W-S-RMM-01", "002010",
    "rv64i_m/F/FCVT-W-S-RNE-01", "002010",
    "rv64i_m/F/FCVT-W-S-RTZ-01", "002010",
    "rv64i_m/F/FCVT-W-S-RUP-01", "002010",
    "rv64i_m/F/FCVT-WU-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FCVT-WU-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FCVT-WU-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FCVT-WU-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FCVT-WU-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FCVT-WU-S-RDN-01", "002010",
    "rv64i_m/F/FCVT-WU-S-RMM-01", "002010",
    "rv64i_m/F/FCVT-WU-S-RNE-01", "002010",
    "rv64i_m/F/FCVT-WU-S-RTZ-01", "002010",
    "rv64i_m/F/FCVT-WU-S-RUP-01", "002010",
    // "rv64i_m/F/FDIV-S-DYN-RDN-01", "002010",
    // "rv64i_m/F/FDIV-S-DYN-RMM-01", "002010",
    // "rv64i_m/F/FDIV-S-DYN-RNE-01", "002010",
    // "rv64i_m/F/FDIV-S-DYN-RTZ-01", "002010",
    // "rv64i_m/F/FDIV-S-DYN-RUP-01", "002010",
    // "rv64i_m/F/FDIV-S-RDN-01", "002010",
    // "rv64i_m/F/FDIV-S-RMM-01", "002010",
    // "rv64i_m/F/FDIV-S-RNE-01", "002010",
    // "rv64i_m/F/FDIV-S-RTZ-01", "002010",
    // "rv64i_m/F/FDIV-S-RUP-01", "002010",
    "rv64i_m/F/FEQ-S-01", "002010",
    "rv64i_m/F/FLE-S-01", "002010",
    "rv64i_m/F/FLT-S-01", "002010",
    "rv64i_m/F/FLW-01", "002210",
    "rv64i_m/F/FMADD-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FMADD-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FMADD-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FMADD-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FMADD-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FMADD-S-RDN-01", "002010",
    "rv64i_m/F/FMADD-S-RMM-01", "002010",
    "rv64i_m/F/FMADD-S-RNE-01", "002010",
    "rv64i_m/F/FMADD-S-RTZ-01", "002010",
    "rv64i_m/F/FMADD-S-RUP-01", "002010",
    "rv64i_m/F/FMAX-S-01", "002010",
    "rv64i_m/F/FMIN-S-01", "002010",
    "rv64i_m/F/FMSUB-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FMSUB-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FMSUB-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FMSUB-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FMSUB-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FMSUB-S-RDN-01", "002010",
    "rv64i_m/F/FMSUB-S-RMM-01", "002010",
    "rv64i_m/F/FMSUB-S-RNE-01", "002010",
    "rv64i_m/F/FMSUB-S-RTZ-01", "002010",
    "rv64i_m/F/FMSUB-S-RUP-01", "002010",
    "rv64i_m/F/FMUL-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FMUL-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FMUL-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FMUL-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FMUL-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FMUL-S-RDN-01", "002010",
    "rv64i_m/F/FMUL-S-RMM-01", "002010",
    "rv64i_m/F/FMUL-S-RNE-01", "002010",
    "rv64i_m/F/FMUL-S-RTZ-01", "002010",
    "rv64i_m/F/FMUL-S-RUP-01", "002010",
    "rv64i_m/F/FMV-W-X-01", "002010",
    "rv64i_m/F/FMV-X-W-01", "002010",
    "rv64i_m/F/FNMADD-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FNMADD-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FNMADD-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FNMADD-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FNMADD-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FNMADD-S-RDN-01", "002010",
    "rv64i_m/F/FNMADD-S-RMM-01", "002010",
    "rv64i_m/F/FNMADD-S-RNE-01", "002010",
    "rv64i_m/F/FNMADD-S-RTZ-01", "002010",
    "rv64i_m/F/FNMADD-S-RUP-01", "002010",
    "rv64i_m/F/FNMSUB-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FNMSUB-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FNMSUB-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FNMSUB-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FNMSUB-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FNMSUB-S-RDN-01", "002010",
    "rv64i_m/F/FNMSUB-S-RMM-01", "002010",
    "rv64i_m/F/FNMSUB-S-RNE-01", "002010",
    "rv64i_m/F/FNMSUB-S-RTZ-01", "002010",
    "rv64i_m/F/FNMSUB-S-RUP-01", "002010",
    "rv64i_m/F/FSGNJN-S-01", "002010",
    "rv64i_m/F/FSGNJ-S-01", "002010",
    "rv64i_m/F/FSGNJX-S-01", "002010",
    // "rv64i_m/F/FSQRT-S-DYN-RDN-01", "002010",
    // "rv64i_m/F/FSQRT-S-DYN-RMM-01", "002010",
    // "rv64i_m/F/FSQRT-S-DYN-RNE-01", "002010",
    // "rv64i_m/F/FSQRT-S-DYN-RTZ-01", "002010",
    // "rv64i_m/F/FSQRT-S-DYN-RUP-01", "002010",
    // "rv64i_m/F/FSQRT-S-RDN-01", "002010",
    // "rv64i_m/F/FSQRT-S-RMM-01", "002010",
    // "rv64i_m/F/FSQRT-S-RNE-01", "002010",
    // "rv64i_m/F/FSQRT-S-RTZ-01", "002010",
    // "rv64i_m/F/FSQRT-S-RUP-01", "002010",
    "rv64i_m/F/FSUB-S-DYN-RDN-01", "002010",
    "rv64i_m/F/FSUB-S-DYN-RMM-01", "002010",
    "rv64i_m/F/FSUB-S-DYN-RNE-01", "002010",
    "rv64i_m/F/FSUB-S-DYN-RTZ-01", "002010",
    "rv64i_m/F/FSUB-S-DYN-RUP-01", "002010",
    "rv64i_m/F/FSUB-S-RDN-01", "002010",
    "rv64i_m/F/FSUB-S-RMM-01", "002010",
    "rv64i_m/F/FSUB-S-RNE-01", "002010",
    "rv64i_m/F/FSUB-S-RTZ-01", "002010",
    "rv64i_m/F/FSUB-S-RUP-01", "002010",
    "rv64i_m/F/FSW-01", "002010"
  };

  string imperas64d[] = '{
    `IMPERASTEST,
    "rv64i_m/D/FADD-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FADD-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FADD-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FADD-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FADD-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FADD-D-RDN-01", "002010",
    "rv64i_m/D/FADD-D-RMM-01", "002010",
    "rv64i_m/D/FADD-D-RNE-01", "002010",
    "rv64i_m/D/FADD-D-RTZ-01", "002010",
    "rv64i_m/D/FADD-D-RUP-01", "002010",
    "rv64i_m/D/FCLASS-D-01", "002010",
    "rv64i_m/D/FCVT-D-L-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-D-L-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-D-L-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-D-L-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-D-L-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-D-L-RDN-01", "002010",
    "rv64i_m/D/FCVT-D-L-RMM-01", "002010",
    "rv64i_m/D/FCVT-D-L-RNE-01", "002010",
    "rv64i_m/D/FCVT-D-L-RTZ-01", "002010",
    "rv64i_m/D/FCVT-D-L-RUP-01", "002010",
    "rv64i_m/D/FCVT-D-LU-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-D-LU-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-D-LU-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-D-LU-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-D-LU-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-D-LU-RDN-01", "002010",
    "rv64i_m/D/FCVT-D-LU-RMM-01", "002010",
    "rv64i_m/D/FCVT-D-LU-RNE-01", "002010",
    "rv64i_m/D/FCVT-D-LU-RTZ-01", "002010",
    "rv64i_m/D/FCVT-D-LU-RUP-01", "002010",
    "rv64i_m/D/FCVT-D-S-01", "002010",
    "rv64i_m/D/FCVT-D-W-01", "002010",
    "rv64i_m/D/FCVT-D-WU-01", "002010",
    "rv64i_m/D/FCVT-L-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-L-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-L-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-L-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-L-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-L-D-RDN-01", "002010",
    "rv64i_m/D/FCVT-L-D-RMM-01", "002010",
    "rv64i_m/D/FCVT-L-D-RNE-01", "002010",
    "rv64i_m/D/FCVT-L-D-RTZ-01", "002010",
    "rv64i_m/D/FCVT-L-D-RUP-01", "002010",
    "rv64i_m/D/FCVT-LU-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-LU-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-LU-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-LU-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-LU-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-LU-D-RDN-01", "002010",
    "rv64i_m/D/FCVT-LU-D-RMM-01", "002010",
    "rv64i_m/D/FCVT-LU-D-RNE-01", "002010",
    "rv64i_m/D/FCVT-LU-D-RTZ-01", "002010",
    "rv64i_m/D/FCVT-LU-D-RUP-01", "002010",
    "rv64i_m/D/FCVT-S-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-S-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-S-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-S-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-S-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-S-D-RDN-01", "002010",
    "rv64i_m/D/FCVT-S-D-RMM-01", "002010",
    "rv64i_m/D/FCVT-S-D-RNE-01", "002010",
    "rv64i_m/D/FCVT-S-D-RTZ-01", "002010",
    "rv64i_m/D/FCVT-S-D-RUP-01", "002010",
    "rv64i_m/D/FCVT-W-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-W-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-W-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-W-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-W-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-W-D-RDN-01", "002010",
    "rv64i_m/D/FCVT-W-D-RMM-01", "002010",
    "rv64i_m/D/FCVT-W-D-RNE-01", "002010",
    "rv64i_m/D/FCVT-W-D-RTZ-01", "002010",
    "rv64i_m/D/FCVT-W-D-RUP-01", "002010",
    "rv64i_m/D/FCVT-WU-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FCVT-WU-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FCVT-WU-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FCVT-WU-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FCVT-WU-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FCVT-WU-D-RDN-01", "002010",
    "rv64i_m/D/FCVT-WU-D-RMM-01", "002010",
    "rv64i_m/D/FCVT-WU-D-RNE-01", "002010",
    "rv64i_m/D/FCVT-WU-D-RTZ-01", "002010",
    "rv64i_m/D/FCVT-WU-D-RUP-01", "002010",
    // "rv64i_m/D/FDIV-D-DYN-RDN-01", "002010",
    // "rv64i_m/D/FDIV-D-DYN-RMM-01", "002010",
    // "rv64i_m/D/FDIV-D-DYN-RNE-01", "002010",
    // "rv64i_m/D/FDIV-D-DYN-RTZ-01", "002010",
    // "rv64i_m/D/FDIV-D-DYN-RUP-01", "002010",
    // "rv64i_m/D/FDIV-D-RDN-01", "002010",
    // "rv64i_m/D/FDIV-D-RMM-01", "002010",
    // "rv64i_m/D/FDIV-D-RNE-01", "002010",
    // "rv64i_m/D/FDIV-D-RTZ-01", "002010",
    // "rv64i_m/D/FDIV-D-RUP-01", "002010",
    "rv64i_m/D/FEQ-D-01", "002010",
    "rv64i_m/D/FLD-01", "002520",
    "rv64i_m/D/FLE-D-01", "002010",
    "rv64i_m/D/FLT-D-01", "002010",
    "rv64i_m/D/FMADD-D-DYN-RDN-01", "003010",
    "rv64i_m/D/FMADD-D-DYN-RMM-01", "003010",
    "rv64i_m/D/FMADD-D-DYN-RNE-01", "003010",
    "rv64i_m/D/FMADD-D-DYN-RTZ-01", "003010",
    "rv64i_m/D/FMADD-D-DYN-RUP-01", "003010",
    "rv64i_m/D/FMADD-D-RDN-01", "003010",
    "rv64i_m/D/FMADD-D-RMM-01", "003010",
    "rv64i_m/D/FMADD-D-RNE-01", "003010",
    "rv64i_m/D/FMADD-D-RTZ-01", "003010",
    "rv64i_m/D/FMADD-D-RUP-01", "003010",
    "rv64i_m/D/FMAX-D-01", "002010",
    "rv64i_m/D/FMIN-D-01", "002010",
    "rv64i_m/D/FMSUB-D-DYN-RDN-01", "003010",
    "rv64i_m/D/FMSUB-D-DYN-RMM-01", "003010",
    "rv64i_m/D/FMSUB-D-DYN-RNE-01", "003010",
    "rv64i_m/D/FMSUB-D-DYN-RTZ-01", "003010",
    "rv64i_m/D/FMSUB-D-DYN-RUP-01", "003010",
    "rv64i_m/D/FMSUB-D-RDN-01", "003010",
    "rv64i_m/D/FMSUB-D-RMM-01", "003010",
    "rv64i_m/D/FMSUB-D-RNE-01", "003010",
    "rv64i_m/D/FMSUB-D-RTZ-01", "003010",
    "rv64i_m/D/FMSUB-D-RUP-01", "003010",
    "rv64i_m/D/FMUL-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FMUL-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FMUL-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FMUL-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FMUL-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FMUL-D-RDN-01", "002010",
    "rv64i_m/D/FMUL-D-RMM-01", "002010",
    "rv64i_m/D/FMUL-D-RNE-01", "002010",
    "rv64i_m/D/FMUL-D-RTZ-01", "002010",
    "rv64i_m/D/FMUL-D-RUP-01", "002010",
    "rv64i_m/D/FMV-D-X-01", "002010",
    "rv64i_m/D/FMV-X-D-01", "002010",
    "rv64i_m/D/FNMADD-D-DYN-RDN-01", "003010",
    "rv64i_m/D/FNMADD-D-DYN-RMM-01", "003010",
    "rv64i_m/D/FNMADD-D-DYN-RNE-01", "003010",
    "rv64i_m/D/FNMADD-D-DYN-RTZ-01", "003010",
    "rv64i_m/D/FNMADD-D-DYN-RUP-01", "003010",
    "rv64i_m/D/FNMADD-D-RDN-01", "003010",
    "rv64i_m/D/FNMADD-D-RMM-01", "003010",
    "rv64i_m/D/FNMADD-D-RNE-01", "003010",
    "rv64i_m/D/FNMADD-D-RTZ-01", "003010",
    "rv64i_m/D/FNMADD-D-RUP-01", "003010",
    "rv64i_m/D/FNMSUB-D-DYN-RDN-01", "003010",
    "rv64i_m/D/FNMSUB-D-DYN-RMM-01", "003010",
    "rv64i_m/D/FNMSUB-D-DYN-RNE-01", "003010",
    "rv64i_m/D/FNMSUB-D-DYN-RTZ-01", "003010",
    "rv64i_m/D/FNMSUB-D-DYN-RUP-01", "003010",
    "rv64i_m/D/FNMSUB-D-RDN-01", "003010",
    "rv64i_m/D/FNMSUB-D-RMM-01", "003010",
    "rv64i_m/D/FNMSUB-D-RNE-01", "003010",
    "rv64i_m/D/FNMSUB-D-RTZ-01", "003010",
    "rv64i_m/D/FNMSUB-D-RUP-01", "003010",
    "rv64i_m/D/FSD-01", "002010",
    "rv64i_m/D/FSGNJ-D-01", "002010",
    "rv64i_m/D/FSGNJN-D-01", "002010",
    "rv64i_m/D/FSGNJX-D-01", "002010",
    // "rv64i_m/D/FSQRT-D-DYN-RDN-01", "002010",
    // "rv64i_m/D/FSQRT-D-DYN-RMM-01", "002010",
    // "rv64i_m/D/FSQRT-D-DYN-RNE-01", "002010",
    // "rv64i_m/D/FSQRT-D-DYN-RTZ-01", "002010",
    // "rv64i_m/D/FSQRT-D-DYN-RUP-01", "002010",
    // "rv64i_m/D/FSQRT-D-RDN-01", "002010",
    // "rv64i_m/D/FSQRT-D-RMM-01", "002010",
    // "rv64i_m/D/FSQRT-D-RNE-01", "002010",
    // "rv64i_m/D/FSQRT-D-RTZ-01", "002010",
    // "rv64i_m/D/FSQRT-D-RUP-01", "002010",
    "rv64i_m/D/FSUB-D-DYN-RDN-01", "002010",
    "rv64i_m/D/FSUB-D-DYN-RMM-01", "002010",
    "rv64i_m/D/FSUB-D-DYN-RNE-01", "002010",
    "rv64i_m/D/FSUB-D-DYN-RTZ-01", "002010",
    "rv64i_m/D/FSUB-D-DYN-RUP-01", "002010",
    "rv64i_m/D/FSUB-D-RDN-01", "002010",
    "rv64i_m/D/FSUB-D-RMM-01", "002010",
    "rv64i_m/D/FSUB-D-RNE-01", "002010",
    "rv64i_m/D/FSUB-D-RTZ-01", "002010",
    "rv64i_m/D/FSUB-D-RUP-01", "002010"
};

  string imperas64m[] = '{
    `IMPERASTEST,
    "rv64i_m/M/DIV-01", "004010",
    "rv64i_m/M/DIVU-01", "004010",
    "rv64i_m/M/DIVUW-01", "003010",
    "rv64i_m/M/DIVW-01", "003010",
    "rv64i_m/M/MUL-01", "004010",
    "rv64i_m/M/MULH-01", "004010",
    "rv64i_m/M/MULHSU-01", "004010",
    "rv64i_m/M/MULHU-01", "004010",
    "rv64i_m/M/MULW-01", "003010",
    "rv64i_m/M/REM-01", "004010",
    "rv64i_m/M/REMU-01", "004010",
    "rv64i_m/M/REMUW-01", "003010",
    "rv64i_m/M/REMW-01", "003010"
  };

  string imperas64c[] = '{
    `IMPERASTEST,
    "rv64i_m/C/C-ADD-01", "003010",
    "rv64i_m/C/C-ADDI-01", "003010",
    "rv64i_m/C/C-ADDI16SP-01", "003010",
    "rv64i_m/C/C-ADDI4SPN-01", "003010",
    "rv64i_m/C/C-ADDIW-01", "003010",
    "rv64i_m/C/C-ADDW-01", "003010",
    "rv64i_m/C/C-AND-01", "003010",
    "rv64i_m/C/C-ANDI-01", "003010",
    "rv64i_m/C/C-BEQZ-01", "004010",
    "rv64i_m/C/C-BNEZ-01", "004010",
    "rv64i_m/C/C-J-01", "003010",
    "rv64i_m/C/C-JALR-01", "004010",
    "rv64i_m/C/C-JR-01", "004010",
    "rv64i_m/C/C-LD-01", "003520",
    "rv64i_m/C/C-LDSP-01", "003520",
    "rv64i_m/C/C-LI-01", "003010",
    "rv64i_m/C/C-LUI-01", "002010",
    "rv64i_m/C/C-LW-01", "003210",
    "rv64i_m/C/C-LWSP-01", "003210",
    "rv64i_m/C/C-MV-01", "003010",
    "rv64i_m/C/C-OR-01", "003010",
    "rv64i_m/C/C-SD-01", "003010",
    "rv64i_m/C/C-SDSP-01", "003010",
    "rv64i_m/C/C-SLLI-01", "003010",
    "rv64i_m/C/C-SRAI-01", "003010",
    "rv64i_m/C/C-SRLI-01", "003010",
    "rv64i_m/C/C-SUB-01", "003010",
    "rv64i_m/C/C-SUBW-01", "003010",
    "rv64i_m/C/C-SW-01", "003010",
    "rv64i_m/C/C-SWSP-01", "003010",
    "rv64i_m/C/C-XOR-01", "003010",
    "rv64i_m/C/I-C-EBREAK-01", "002000",
    "rv64i_m/C/I-C-NOP-01", "002000"
  };

  string imperas64iNOc[] = {
    `IMPERASTEST,
    "rv64i_m/I/I-MISALIGN_JMP-01", "002000"
  };

  string imperas64i[] = '{
    `IMPERASTEST,
    "rv64i_m/I/I-DELAY_SLOTS-01", "002010",
    "rv64i_m/I/ADD-01", "004010",
    "rv64i_m/I/ADDI-01", "003010",
    "rv64i_m/I/ADDIW-01", "003010",
    "rv64i_m/I/ADDW-01", "003010",
    "rv64i_m/I/AND-01", "004010",
    "rv64i_m/I/ANDI-01", "003010",
    "rv64i_m/I/AUIPC-01", "003010",
    "rv64i_m/I/BEQ-01", "005010",
    "rv64i_m/I/BGE-01", "005010",
    "rv64i_m/I/BGEU-01", "005010",
    "rv64i_m/I/BLT-01", "005010",
    "rv64i_m/I/BLTU-01", "005010",
    "rv64i_m/I/BNE-01", "005010",
    "rv64i_m/I/I-DELAY_SLOTS-01", "002010",
    "rv64i_m/I/I-EBREAK-01", "002010",
    "rv64i_m/I/I-ECALL-01", "002010",
    "rv64i_m/I/I-ENDIANESS-01", "002010",
    "rv64i_m/I/I-IO-01", "002050",
//    "rv64i_m/I/I-MISALIGN_JMP-01", "002000",
    "rv64i_m/I/I-MISALIGN_LDST-01", "002010",
    "rv64i_m/I/I-NOP-01", "002000",
    "rv64i_m/I/I-RF_size-01", "002000",
    "rv64i_m/I/I-RF_width-01", "002000",
    "rv64i_m/I/I-RF_x0-01", "002010",
    "rv64i_m/I/JAL-01", "004010",
    "rv64i_m/I/JALR-01", "005010",
    "rv64i_m/I/LB-01", "004120",
    "rv64i_m/I/LBU-01", "004120",
    "rv64i_m/I/LD-01", "004520",
    "rv64i_m/I/LH-01", "004150",
    "rv64i_m/I/LHU-01", "004150",
    "rv64i_m/I/LUI-01", "002010",
    "rv64i_m/I/LW-01", "004210",
    "rv64i_m/I/LWU-01", "004210",
    "rv64i_m/I/OR-01", "004010",
    "rv64i_m/I/ORI-01", "003010",
    "rv64i_m/I/SB-01", "004010",
    "rv64i_m/I/SD-01", "004010",
    "rv64i_m/I/SH-01", "004010",
    "rv64i_m/I/SLL-01", "003010",
    "rv64i_m/I/SLLI-01", "003010",
    "rv64i_m/I/SLLIW-01", "003010",
    "rv64i_m/I/SLLW-01", "003010",
    "rv64i_m/I/SLT-01", "004010",
    "rv64i_m/I/SLTI-01", "003010",
    "rv64i_m/I/SLTIU-01", "003010",
    "rv64i_m/I/SLTU-01", "004010",
    "rv64i_m/I/SRA-01", "003010",
    "rv64i_m/I/SRAI-01", "003010",
    "rv64i_m/I/SRAIW-01", "003010",
    "rv64i_m/I/SRAW-01", "003010",
    "rv64i_m/I/SRL-01", "003010",
    "rv64i_m/I/SRLI-01", "003010",
    "rv64i_m/I/SRLIW-01", "003010",
    "rv64i_m/I/SRLW-01", "003010",
    "rv64i_m/I/SUB-01", "004010",
    "rv64i_m/I/SUBW-01", "003010",
    "rv64i_m/I/SW-01", "004010",
    "rv64i_m/I/XOR-01", "004010",
    "rv64i_m/I/XORI-01", "003010"
  };

  string imperas32m[] = '{
    `IMPERASTEST,
    "rv32i_m/M/DIV-01", "002010",
    "rv32i_m/M/DIVU-01", "002010",
    "rv32i_m/M/MUL-01", "002010",
    "rv32i_m/M/MULH-01", "002010",
    "rv32i_m/M/MULHSU-01", "002010",
    "rv32i_m/M/MULHU-01", "002010",
    "rv32i_m/M/REM-01", "002010",
    "rv32i_m/M/REMU-01", "002010"
  };

  string imperas32c[] = '{
    `IMPERASTEST,
    "rv32i_m/C/C-ADD-01", "002010",
    "rv32i_m/C/C-ADDI-01", "002010",
    "rv32i_m/C/C-ADDI16SP-01", "002010",
    "rv32i_m/C/C-ADDI4SPN-01", "002010",
    "rv32i_m/C/C-AND-01", "002010",
    "rv32i_m/C/C-ANDI-01", "002010",
    "rv32i_m/C/C-BEQZ-01", "003010",
    "rv32i_m/C/C-BNEZ-01", "003010",
    "rv32i_m/C/C-J-01", "002010",
    "rv32i_m/C/C-JAL-01", "002010",
    "rv32i_m/C/C-JALR-01", "003010",
    "rv32i_m/C/C-JR-01", "003010",
    "rv32i_m/C/C-LI-01", "002010",
    "rv32i_m/C/C-LUI-01", "002010",
    "rv32i_m/C/C-LW-01", "002120",
    "rv32i_m/C/C-LWSP-01", "002120",
    "rv32i_m/C/C-MV-01", "002010",
    "rv32i_m/C/C-OR-01", "002010",
    "rv32i_m/C/C-SLLI-01", "002010",
    "rv32i_m/C/C-SRAI-01", "002010",
    "rv32i_m/C/C-SRLI-01", "002010",
    "rv32i_m/C/C-SUB-01", "002010",
    "rv32i_m/C/C-SW-01", "002010",
    "rv32i_m/C/C-SWSP-01", "002010",
    "rv32i_m/C/C-XOR-01", "002010",
    "rv32i_m/C/I-C-EBREAK-01", "002000",
    "rv32i_m/C/I-C-NOP-01", "002000"
  };

  string imperas32iNOc[] = {
    `IMPERASTEST,
    "rv32i_m/I/I-MISALIGN_JMP-01", "002000"
  };

  string imperas32i[] = {
    `IMPERASTEST,
    "rv32i_m/I/ADD-01", "002010",
    "rv32i_m/I/ADDI-01", "002010",
    "rv32i_m/I/AND-01", "002010",
    "rv32i_m/I/ANDI-01", "002010",
    "rv32i_m/I/AUIPC-01", "002010",
    "rv32i_m/I/BEQ-01", "003010",
    "rv32i_m/I/BGE-01", "003010",
    "rv32i_m/I/BGEU-01", "003010",
    "rv32i_m/I/BLT-01", "003010",
    "rv32i_m/I/BLTU-01", "003010",
    "rv32i_m/I/BNE-01", "003010",
    "rv32i_m/I/I-DELAY_SLOTS-01", "002010",
    "rv32i_m/I/I-EBREAK-01", "002010",
    "rv32i_m/I/I-ECALL-01", "002010",
    "rv32i_m/I/I-ENDIANESS-01", "002010",
    "rv32i_m/I/I-IO-01", "002030",
//    "rv32i_m/I/I-MISALIGN_JMP-01", "002000",
    "rv32i_m/I/I-MISALIGN_LDST-01", "002010",
    "rv32i_m/I/I-NOP-01", "002000",
    "rv32i_m/I/I-RF_size-01", "002000",
    "rv32i_m/I/I-RF_width-01", "002000",
    "rv32i_m/I/I-RF_x0-01", "002010",
    "rv32i_m/I/JAL-01", "003010",
    "rv32i_m/I/JALR-01", "003010",
    "rv32i_m/I/LB-01", "003030",
    "rv32i_m/I/LBU-01", "003030",
    "rv32i_m/I/LH-01", "003060",
    "rv32i_m/I/LHU-01", "003060",
    "rv32i_m/I/LUI-01", "002010",
    "rv32i_m/I/LW-01", "003120",
    "rv32i_m/I/OR-01", "002010",
    "rv32i_m/I/ORI-01", "002010",
    "rv32i_m/I/SB-01", "003010",
    "rv32i_m/I/SH-01", "003010",
    "rv32i_m/I/SLL-01", "002010",
    "rv32i_m/I/SLLI-01", "002010",
    "rv32i_m/I/SLT-01", "002010",
    "rv32i_m/I/SLTI-01", "002010",
    "rv32i_m/I/SLTIU-01", "002010",
    "rv32i_m/I/SLTU-01", "002010",
    "rv32i_m/I/SRA-01", "002010",
    "rv32i_m/I/SRAI-01", "002010",
    "rv32i_m/I/SRL-01", "002010",
    "rv32i_m/I/SRLI-01", "002010",
    "rv32i_m/I/SUB-01", "002010",
    "rv32i_m/I/SW-01", "003010",
    "rv32i_m/I/XOR-01", "002010",
    "rv32i_m/I/XORI-01", "002010"   
  };

  string testsBP64[] = '{
    `IMPERASTEST,
    "rv64BP/simple", "10000",
    "rv64BP/mmm", "1000000",
    "rv64BP/linpack_bench", "1000000",
    "rv64BP/sieve", "1000000",
    "rv64BP/qsort", "1000000",
    "rv64BP/dhrystone", "1000000"
  };

  string imperas32p[] = '{
    `MYIMPERASTEST,
    "rv32p/WALLY-MSTATUS", "2000",
    "rv32p/WALLY-MCAUSE", "3000",
    "rv32p/WALLY-SCAUSE", "2000",
    "rv32p/WALLY-MEPC", "5000",
    "rv32p/WALLY-SEPC", "4000",
    "rv32p/WALLY-MTVAL", "5000",
    "rv32p/WALLY-STVAL", "4000",
    "rv32p/WALLY-MARCHID", "4000",
    "rv32p/WALLY-MIMPID", "4000",
    "rv32p/WALLY-MHARTID", "4000",
    "rv32p/WALLY-MVENDORID", "4000",
    "rv32p/WALLY-MTVEC", "2000",
    "rv32p/WALLY-STVEC", "2000",
    "rv32p/WALLY-MIE", "3000",
    "rv32p/WALLY-MEDELEG", "4000",
    "rv32p/WALLY-IP", "3000",
    "rv32p/WALLY-CSR-PERMISSIONS-M", "5000",
    "rv32p/WALLY-CSR-PERMISSIONS-S", "3000"
  };

  string arch64priv[] = '{
    `RISCVARCHTEST,
    "rv64i_m/privilege/ebreak", "2090",
    "rv64i_m/privilege/ecall", "2090",
    "rv64i_m/privilege/misalign-beq-01", "20a0",
    "rv64i_m/privilege/misalign-bge-01", "20a0",
    "rv64i_m/privilege/misalign-bgeu-01", "20a0",
    "rv64i_m/privilege/misalign-blt-01", "20a0",
    "rv64i_m/privilege/misalign-bltu-01", "20a0",
    "rv64i_m/privilege/misalign-bne-01", "20a0",
    "rv64i_m/privilege/misalign-jal-01", "20a0",
    "rv64i_m/privilege/misalign-ld-01", "20a0",
    "rv64i_m/privilege/misalign-lh-01", "20a0",
    "rv64i_m/privilege/misalign-lhu-01", "20a0",
    "rv64i_m/privilege/misalign-lw-01", "20a0",
    "rv64i_m/privilege/misalign-lwu-01", "20a0",
    "rv64i_m/privilege/misalign-sd-01", "20a0",
    "rv64i_m/privilege/misalign-sh-01", "20a0",
    "rv64i_m/privilege/misalign-sw-01", "20a0",
    "rv64i_m/privilege/misalign1-jalr-01", "20a0",
    "rv64i_m/privilege/misalign2-jalr-01", "20a0"
    };

  string arch64m[] = '{
    `RISCVARCHTEST,
    "rv64i_m/M/div-01", "9010",
    "rv64i_m/M/divu-01", "a010",
    "rv64i_m/M/divuw-01", "a010",
    "rv64i_m/M/divw-01", "9010",
    "rv64i_m/M/mul-01", "9010",
    "rv64i_m/M/mulh-01", "9010",
    "rv64i_m/M/mulhsu-01", "9010",
    "rv64i_m/M/mulhu-01", "a010",
    "rv64i_m/M/mulw-01", "9010",
    "rv64i_m/M/rem-01", "9010",
    "rv64i_m/M/remu-01", "a010",
    "rv64i_m/M/remuw-01", "a010",
    "rv64i_m/M/remw-01", "9010"
   };

  string arch64c[] = '{
    `RISCVARCHTEST,
    "rv64i_m/C/cadd-01", "8010",
    "rv64i_m/C/caddi-01", "4010",
    "rv64i_m/C/caddi16sp-01", "2010",
    "rv64i_m/C/caddi4spn-01", "2010",
    "rv64i_m/C/caddiw-01", "4010",
    "rv64i_m/C/caddw-01", "8010",
    "rv64i_m/C/cand-01", "8010",
    "rv64i_m/C/candi-01", "4010",
    "rv64i_m/C/cbeqz-01", "4010",
    "rv64i_m/C/cbnez-01", "5010",
    "rv64i_m/C/cj-01", "3010",
    "rv64i_m/C/cjalr-01", "2010",
    "rv64i_m/C/cjr-01", "2010",
    "rv64i_m/C/cld-01", "2010",
    "rv64i_m/C/cldsp-01", "2010",
    "rv64i_m/C/cli-01", "2010",
    "rv64i_m/C/clui-01", "2010",
    "rv64i_m/C/clw-01", "2010",
    "rv64i_m/C/clwsp-01", "2010",
    "rv64i_m/C/cmv-01", "2010",
    "rv64i_m/C/cnop-01", "2010",
    "rv64i_m/C/cor-01", "8010",
    "rv64i_m/C/csd-01", "3010",
    "rv64i_m/C/csdsp-01", "3010",
    "rv64i_m/C/cslli-01", "2010",
    "rv64i_m/C/csrai-01", "2010",
    "rv64i_m/C/csrli-01", "2010",
    "rv64i_m/C/csub-01", "8010",
    "rv64i_m/C/csubw-01", "8010",
    "rv64i_m/C/csw-01", "3010",
    "rv64i_m/C/cswsp-01", "3010",
    "rv64i_m/C/cxor-01", "8010"
  };

  string arch64cpriv[] = '{
//    `RISCVARCHTEST,
      "rv64i_m/C/cebreak-01", "2070"
  };

  string arch64i[] = '{
    `RISCVARCHTEST,
    "rv64i_m/I/add-01", "9010",
    "rv64i_m/I/addi-01", "6010",
    "rv64i_m/I/addiw-01", "6010",
    "rv64i_m/I/addw-01", "9010",
    "rv64i_m/I/and-01", "9010",
    "rv64i_m/I/andi-01", "6010",
    "rv64i_m/I/auipc-01", "2010",
    "rv64i_m/I/beq-01", "47010",
    "rv64i_m/I/bge-01", "46010",
    "rv64i_m/I/bgeu-01", "56010",
    "rv64i_m/I/blt-01", "4d010",
    "rv64i_m/I/bltu-01", "57010",
    "rv64i_m/I/bne-01", "43010",
    "rv64i_m/I/fence-01", "2010",
    "rv64i_m/I/jal-01", "122010",
    "rv64i_m/I/jalr-01", "2010",
    "rv64i_m/I/lb-align-01", "2010",
    "rv64i_m/I/lbu-align-01", "2010",
    "rv64i_m/I/ld-align-01", "2010",
    "rv64i_m/I/lh-align-01", "2010",
    "rv64i_m/I/lhu-align-01", "2010",
    "rv64i_m/I/lui-01", "2010",
    "rv64i_m/I/lw-align-01", "2010",
    "rv64i_m/I/lwu-align-01", "2010",
    "rv64i_m/I/or-01", "9010",
    "rv64i_m/I/ori-01", "6010",
    "rv64i_m/I/sb-align-01", "3010",
    "rv64i_m/I/sd-align-01", "3010",
    "rv64i_m/I/sh-align-01", "3010",
    "rv64i_m/I/sll-01", "3010",
    "rv64i_m/I/slli-01", "2010",
    "rv64i_m/I/slliw-01", "2010",
    "rv64i_m/I/sllw-01", "3010",
    "rv64i_m/I/slt-01", "9010",
    "rv64i_m/I/slti-01", "6010",
    "rv64i_m/I/sltiu-01", "6010",
    "rv64i_m/I/sltu-01", "a010",
    "rv64i_m/I/sra-01", "3010",
    "rv64i_m/I/srai-01", "2010",
    "rv64i_m/I/sraiw-01", "2010",
    "rv64i_m/I/sraw-01", "3010",
    "rv64i_m/I/srl-01", "3010",
    "rv64i_m/I/srli-01", "2010",
    "rv64i_m/I/srliw-01", "2010",
    "rv64i_m/I/srlw-01", "3010",
    "rv64i_m/I/sub-01", "9010",
    "rv64i_m/I/subw-01", "9010",
    "rv64i_m/I/sw-align-01", "3010",
    "rv64i_m/I/xor-01", "9010",
    "rv64i_m/I/xori-01", "6010"
  };


  string arch64d[] = '{
    `RISCVARCHTEST,
    "rv64i_m/D/d_fadd_b10-01", "8690",
    "rv64i_m/D/d_fadd_b1-01", "8430",
    "rv64i_m/D/d_fadd_b11-01", "74da0", 
    "rv64i_m/D/d_fadd_b12-01", "2350",
    "rv64i_m/D/d_fadd_b13-01", "3cb0",
    "rv64i_m/D/d_fadd_b2-01", "5160",
    "rv64i_m/D/d_fadd_b3-01", "d640",
    "rv64i_m/D/d_fadd_b4-01", "3900",
    "rv64i_m/D/d_fadd_b5-01", "3d50",
    "rv64i_m/D/d_fadd_b7-01", "5530",
    "rv64i_m/D/d_fadd_b8-01", "11c10",
    "rv64i_m/D/d_fclass_b1-01", "2110",
    "rv64i_m/D/d_fcvt.d.l_b25-01", "2110",
    "rv64i_m/D/d_fcvt.d.l_b26-01", "2220",
    "rv64i_m/D/d_fcvt.d.lu_b25-01", "2110",
    "rv64i_m/D/d_fcvt.d.lu_b26-01", "2220",
    "rv64i_m/D/d_fcvt.d.s_b1-01", "2110", 
    "rv64i_m/D/d_fcvt.d.s_b22-01", "2110", 
    "rv64i_m/D/d_fcvt.d.s_b23-01", "2110",
    "rv64i_m/D/d_fcvt.d.s_b24-01", "2110",
    "rv64i_m/D/d_fcvt.d.s_b27-01", "2110",
    "rv64i_m/D/d_fcvt.d.s_b28-01", "2110",
    "rv64i_m/D/d_fcvt.d.s_b29-01", "2110", 
    "rv64i_m/D/d_fcvt.d.w_b25-01", "2120",
    "rv64i_m/D/d_fcvt.d.w_b26-01", "2220",
    "rv64i_m/D/d_fcvt.d.wu_b25-01", "2110",
    "rv64i_m/D/d_fcvt.d.wu_b26-01", "2220", 
    "rv64i_m/D/d_fcvt.l.d_b1-01", "2120",
    "rv64i_m/D/d_fcvt.l.d_b22-01", "2260",
    "rv64i_m/D/d_fcvt.l.d_b23-01", "2180",
    "rv64i_m/D/d_fcvt.l.d_b24-01", "2360", 
    "rv64i_m/D/d_fcvt.l.d_b27-01", "2110",
    "rv64i_m/D/d_fcvt.l.d_b28-01", "2120",
    "rv64i_m/D/d_fcvt.l.d_b29-01", "22a0",
    "rv64i_m/D/d_fcvt.lu.d_b1-01", "2120", 
    "rv64i_m/D/d_fcvt.lu.d_b22-01", "2260",
    "rv64i_m/D/d_fcvt.lu.d_b23-01", "2180",
    "rv64i_m/D/d_fcvt.lu.d_b24-01", "2360", 
    "rv64i_m/D/d_fcvt.lu.d_b27-01", "2120",
    "rv64i_m/D/d_fcvt.lu.d_b28-01", "2120",
    "rv64i_m/D/d_fcvt.lu.d_b29-01", "22a0",
    "rv64i_m/D/d_fcvt.s.d_b1-01", "2110",
    "rv64i_m/D/d_fcvt.s.d_b22-01", "2110",
    "rv64i_m/D/d_fcvt.s.d_b23-01", "2180",
    "rv64i_m/D/d_fcvt.s.d_b24-01", "2360",
    "rv64i_m/D/d_fcvt.s.d_b27-01", "2110",
    "rv64i_m/D/d_fcvt.s.d_b28-01", "2110",
    "rv64i_m/D/d_fcvt.s.d_b29-01", "22a0",
    "rv64i_m/D/d_fcvt.w.d_b1-01", "2120", 
    "rv64i_m/D/d_fcvt.w.d_b22-01", "2160", 
    "rv64i_m/D/d_fcvt.w.d_b23-01", "2180",
    "rv64i_m/D/d_fcvt.w.d_b24-01", "2360",
    "rv64i_m/D/d_fcvt.w.d_b27-01", "2120",
    "rv64i_m/D/d_fcvt.w.d_b28-01", "2120",
    "rv64i_m/D/d_fcvt.w.d_b29-01", "22a0",
    "rv64i_m/D/d_fcvt.wu.d_b1-01", "2120", 
    "rv64i_m/D/d_fcvt.wu.d_b22-01", "2160",
    "rv64i_m/D/d_fcvt.wu.d_b23-01", "2180",
    "rv64i_m/D/d_fcvt.wu.d_b24-01", "2360", 
    "rv64i_m/D/d_fcvt.wu.d_b27-01", "2120",
    "rv64i_m/D/d_fcvt.wu.d_b28-01", "2120",
    "rv64i_m/D/d_fcvt.wu.d_b29-01", "22a0",
    // "rv64i_m/D/d_fdiv_b1-01", "8430", // RV NaNs need to be positive
    // "rv64i_m/D/d_fdiv_b20-01", "3fa0", // looks like flags
    // "rv64i_m/D/d_fdiv_b2-01", "5170", // also flags
    // "rv64i_m/D/d_fdiv_b21-01", "8a70", // positive NaNs again
    "rv64i_m/D/d_fdiv_b3-01", "d630",
    // "rv64i_m/D/d_fdiv_b4-01", "38f0", // flags
    "rv64i_m/D/d_fdiv_b5-01", "3d50",
    // "rv64i_m/D/d_fdiv_b6-01", "38f0", // flags
    "rv64i_m/D/d_fdiv_b7-01", "5530",
    // "rv64i_m/D/d_fdiv_b8-01", "11c10", // flags
    // "rv64i_m/D/d_fdiv_b9-01", "1b0f0",  might be a flag too
    "rv64i_m/D/d_feq_b1-01", "7430",
    "rv64i_m/D/d_feq_b19-01", "c4c0",
    "rv64i_m/D/d_fld-align-01", "2010",
    "rv64i_m/D/d_fle_b1-01", "7430",
    "rv64i_m/D/d_fle_b19-01", "c4c0",
    "rv64i_m/D/d_flt_b1-01", "7430",
    "rv64i_m/D/d_flt_b19-01", "d800",
    "rv64i_m/D/d_fmadd_b14-01", "3fd0",
    "rv64i_m/D/d_fmadd_b16-01", "43b0",
    "rv64i_m/D/d_fmadd_b17-01", "43b0", 
    "rv64i_m/D/d_fmadd_b18-01", "5a20", 
    "rv64i_m/D/d_fmadd_b2-01", "5ab0",
    "rv64i_m/D/d_fmadd_b3-01", "119d0",
    "rv64i_m/D/d_fmadd_b4-01", "3df0",
    "rv64i_m/D/d_fmadd_b5-01", "4480",
    "rv64i_m/D/d_fmadd_b6-01", "3df0",
    "rv64i_m/D/d_fmadd_b7-01", "6050",
    "rv64i_m/D/d_fmadd_b8-01", "15aa0",
    "rv64i_m/D/d_fmax_b1-01", "8430",
    "rv64i_m/D/d_fmax_b19-01", "d5c0",
    "rv64i_m/D/d_fmin_b1-01", "8430",
    "rv64i_m/D/d_fmin_b19-01", "d4b0",
    "rv64i_m/D/d_fmsub_b14-01", "3fd0",
    "rv64i_m/D/d_fmsub_b16-01", "43b0", 
    "rv64i_m/D/d_fmsub_b17-01", "43b0",
    "rv64i_m/D/d_fmsub_b18-01", "5a20", 
    "rv64i_m/D/d_fmsub_b2-01", "5ab0",
    "rv64i_m/D/d_fmsub_b3-01", "119f0",
    "rv64i_m/D/d_fmsub_b4-01", "3df0",
    "rv64i_m/D/d_fmsub_b5-01", "4480",
    "rv64i_m/D/d_fmsub_b6-01", "3df0",
    "rv64i_m/D/d_fmsub_b7-01", "6050",
    "rv64i_m/D/d_fmsub_b8-01", "15aa0",
    "rv64i_m/D/d_fmul_b1-01", "8430",
    "rv64i_m/D/d_fmul_b2-01", "5180",
    "rv64i_m/D/d_fmul_b3-01", "d640",
    "rv64i_m/D/d_fmul_b4-01", "38f0",
    "rv64i_m/D/d_fmul_b5-01", "3d50",
    "rv64i_m/D/d_fmul_b6-01", "38f0",
    "rv64i_m/D/d_fmul_b7-01", "5540",
    "rv64i_m/D/d_fmul_b8-01", "11c10",
    "rv64i_m/D/d_fmul_b9-01", "1b0f0",
    "rv64i_m/D/d_fmv.d.x_b25-01", "2110",
    "rv64i_m/D/d_fmv.d.x_b26-01", "2220",
    "rv64i_m/D/d_fmv.x.d_b1-01", "2120",
    "rv64i_m/D/d_fmv.x.d_b22-01", "2110",
    "rv64i_m/D/d_fmv.x.d_b23-01", "2110",
    "rv64i_m/D/d_fmv.x.d_b24-01", "2120",
    "rv64i_m/D/d_fmv.x.d_b27-01", "2120",
    "rv64i_m/D/d_fmv.x.d_b28-01", "2110",
    "rv64i_m/D/d_fmv.x.d_b29-01", "2120",
    "rv64i_m/D/d_fnmadd_b14-01", "3fd0",
    "rv64i_m/D/d_fnmadd_b16-01", "4390",
    "rv64i_m/D/d_fnmadd_b17-01", "4390",
    "rv64i_m/D/d_fnmadd_b18-01", "5a20", 
    "rv64i_m/D/d_fnmadd_b2-01", "5ab0",
    "rv64i_m/D/d_fnmadd_b3-01", "119d0", 
    "rv64i_m/D/d_fnmadd_b4-01", "3df0",
    "rv64i_m/D/d_fnmadd_b5-01", "4480",
    "rv64i_m/D/d_fnmadd_b6-01", "3df0",
    "rv64i_m/D/d_fnmadd_b7-01", "6050",
    "rv64i_m/D/d_fnmadd_b8-01", "15aa0",
    "rv64i_m/D/d_fnmsub_b14-01", "3fd0",
    "rv64i_m/D/d_fnmsub_b16-01", "4390",
    "rv64i_m/D/d_fnmsub_b17-01", "4390", 
    "rv64i_m/D/d_fnmsub_b18-01", "5a20",
    "rv64i_m/D/d_fnmsub_b2-01", "5aa0",
    "rv64i_m/D/d_fnmsub_b3-01", "119d0",
    "rv64i_m/D/d_fnmsub_b4-01", "3e20",
    "rv64i_m/D/d_fnmsub_b5-01", "4480",
    "rv64i_m/D/d_fnmsub_b6-01", "3e10",
    "rv64i_m/D/d_fnmsub_b7-01", "6050",
    "rv64i_m/D/d_fnmsub_b8-01", "15aa0", 
    "rv64i_m/D/d_fsd-align-01", "2010",
    "rv64i_m/D/d_fsgnj_b1-01", "8430",
    "rv64i_m/D/d_fsgnjn_b1-01", "8430",
    "rv64i_m/D/d_fsgnjx_b1-01", "8430",
    // "rv64i_m/D/d_fsqrt_b1-01", "2110", // flg
    // "rv64i_m/D/d_fsqrt_b20-01", "3460", // flg
    // "rv64i_m/D/d_fsqrt_b2-01", "2190", // flg - I'm going to stop here with the sqrt
    // "rv64i_m/D/d_fsqrt_b3-01", "2120",
    // "rv64i_m/D/d_fsqrt_b4-01", "2110",
    // "rv64i_m/D/d_fsqrt_b5-01", "2110",
    // "rv64i_m/D/d_fsqrt_b7-01", "2110",
    // "rv64i_m/D/d_fsqrt_b8-01", "2110",
    // "rv64i_m/D/d_fsqrt_b9-01", "4c10",
    "rv64i_m/D/d_fsub_b10-01", "8660",
    "rv64i_m/D/d_fsub_b1-01", "8440",
    "rv64i_m/D/d_fsub_b11-01", "74da0",
    "rv64i_m/D/d_fsub_b12-01", "2350",
    "rv64i_m/D/d_fsub_b13-01", "3cb0",
    "rv64i_m/D/d_fsub_b2-01", "5160",
    "rv64i_m/D/d_fsub_b3-01", "d630",
    "rv64i_m/D/d_fsub_b4-01", "38f0",
    "rv64i_m/D/d_fsub_b5-01", "3d50",
    "rv64i_m/D/d_fsub_b7-01", "5530",
    "rv64i_m/D/d_fsub_b8-01", "11c10"
  };

    string arch32priv[] = '{
    `RISCVARCHTEST,
    "rv32i_m/privilege/ebreak", "2070",
    "rv32i_m/privilege/ecall", "2070",
    "rv32i_m/privilege/misalign-beq-01", "2080",
    "rv32i_m/privilege/misalign-bge-01", "2080",
    "rv32i_m/privilege/misalign-bgeu-01", "2080",
    "rv32i_m/privilege/misalign-blt-01", "2080",
    "rv32i_m/privilege/misalign-bltu-01", "2080",
    "rv32i_m/privilege/misalign-bne-01", "2080",
    "rv32i_m/privilege/misalign-jal-01", "2080",
    "rv32i_m/privilege/misalign-lh-01", "2080",
    "rv32i_m/privilege/misalign-lhu-01", "2080",
    "rv32i_m/privilege/misalign-lw-01", "2080",
    "rv32i_m/privilege/misalign-sh-01", "2080",
    "rv32i_m/privilege/misalign-sw-01", "2080",
    "rv32i_m/privilege/misalign1-jalr-01", "2080",
    "rv32i_m/privilege/misalign2-jalr-01", "2080"
    };

  string arch32m[] = '{
    `RISCVARCHTEST,
    "rv32i_m/M/div-01", "5010",
    "rv32i_m/M/divu-01", "5010",
    "rv32i_m/M/mul-01", "5010",
    "rv32i_m/M/mulh-01", "5010",
    "rv32i_m/M/mulhsu-01", "5010",
    "rv32i_m/M/mulhu-01", "5010",
    "rv32i_m/M/rem-01", "5010",
    "rv32i_m/M/remu-01", "5010"
   };

  string arch32f[] = '{
    `RISCVARCHTEST,
    "rv32i_m/F/fadd_b1-01", "7220",
    "rv32i_m/F/fadd_b10-01", "2270", 
    "rv32i_m/F/fadd_b11-01", "3fb40",
    "rv32i_m/F/fadd_b12-01", "21b0",
    "rv32i_m/F/fadd_b13-01", "3660",
    "rv32i_m/F/fadd_b2-01", "38b0",
    "rv32i_m/F/fadd_b3-01", "b320",
    "rv32i_m/F/fadd_b4-01", "3480",
    "rv32i_m/F/fadd_b5-01", "3700",
    "rv32i_m/F/fadd_b7-01", "3520",
    "rv32i_m/F/fadd_b8-01", "104a0",
    "rv32i_m/F/fclass_b1-01", "2090",
    "rv32i_m/F/fcvt.s.w_b25-01", "20a0",
    "rv32i_m/F/fcvt.s.w_b26-01", "3290",
    "rv32i_m/F/fcvt.s.wu_b25-01", "20a0",
    "rv32i_m/F/fcvt.s.wu_b26-01", "3290",
    "rv32i_m/F/fcvt.w.s_b1-01", "2090",
    "rv32i_m/F/fcvt.w.s_b22-01", "20b0",
    "rv32i_m/F/fcvt.w.s_b23-01", "20c0",
    "rv32i_m/F/fcvt.w.s_b24-01", "21b0",
    "rv32i_m/F/fcvt.w.s_b27-01", "2090",
    "rv32i_m/F/fcvt.w.s_b28-01", "2090",
    "rv32i_m/F/fcvt.w.s_b29-01", "2150",
    "rv32i_m/F/fcvt.wu.s_b1-01", "2090",
    "rv32i_m/F/fcvt.wu.s_b22-01", "20b0",
    "rv32i_m/F/fcvt.wu.s_b23-01", "20c0",
    "rv32i_m/F/fcvt.wu.s_b24-01", "21b0",
    "rv32i_m/F/fcvt.wu.s_b27-01", "2090",
    "rv32i_m/F/fcvt.wu.s_b28-01", "2090",
    "rv32i_m/F/fcvt.wu.s_b29-01", "2150",
    // "rv32i_m/F/fdiv_b1-01", "7220", // NaN i'm going to skip div, probably the same problems as the double version
    // "rv32i_m/F/fdiv_b2-01", "2350",
    // "rv32i_m/F/fdiv_b20-01", "38c0",
    // "rv32i_m/F/fdiv_b21-01", "7540",
    // "rv32i_m/F/fdiv_b3-01", "b320",
    // "rv32i_m/F/fdiv_b4-01", "3480",
    // "rv32i_m/F/fdiv_b5-01", "3700",
    // "rv32i_m/F/fdiv_b6-01", "3480",
    // "rv32i_m/F/fdiv_b7-01", "3520",
    // "rv32i_m/F/fdiv_b8-01", "104a0",
    // "rv32i_m/F/fdiv_b9-01", "d960",
    "rv32i_m/F/feq_b1-01", "6220",
    "rv32i_m/F/feq_b19-01", "a190",
    "rv32i_m/F/fle_b1-01", "6220",
    "rv32i_m/F/fle_b19-01", "a190",
    "rv32i_m/F/flt_b1-01", "6220",
    "rv32i_m/F/flt_b19-01", "8ee0", 
    "rv32i_m/F/flw-align-01", "2010",
    "rv32i_m/F/fmadd_b1-01", "96860",
    "rv32i_m/F/fmadd_b14-01", "23d0",
// --passes but is timeconsuming    "rv32i_m/F/fmadd_b15-01", "19bb30",
    "rv32i_m/F/fmadd_b16-01", "39d0",
    "rv32i_m/F/fmadd_b17-01", "39d0",
    "rv32i_m/F/fmadd_b18-01", "4d10", 
    "rv32i_m/F/fmadd_b2-01", "4d60",
    "rv32i_m/F/fmadd_b3-01", "d4f0",
    "rv32i_m/F/fmadd_b4-01", "3700",
    "rv32i_m/F/fmadd_b5-01", "3ac0",
    "rv32i_m/F/fmadd_b6-01", "3700",
    "rv32i_m/F/fmadd_b7-01", "37f0",
    "rv32i_m/F/fmadd_b8-01", "13f30", 
    "rv32i_m/F/fmax_b1-01", "7220",
    "rv32i_m/F/fmax_b19-01", "9e00",
    "rv32i_m/F/fmin_b1-01", "7220",
    "rv32i_m/F/fmin_b19-01", "9f20",
    "rv32i_m/F/fmsub_b1-01", "96860",
    "rv32i_m/F/fmsub_b14-01", "23d0",
    "rv32i_m/F/fmsub_b15-01", "19bb30",
    "rv32i_m/F/fmsub_b16-01", "39d0",
    "rv32i_m/F/fmsub_b17-01", "39d0",
    "rv32i_m/F/fmsub_b18-01", "4d20", 
    "rv32i_m/F/fmsub_b2-01", "4d60",
    "rv32i_m/F/fmsub_b3-01", "d4f0",
    "rv32i_m/F/fmsub_b4-01", "3700",
    "rv32i_m/F/fmsub_b5-01", "3ac0",
    "rv32i_m/F/fmsub_b6-01", "3700", 
    "rv32i_m/F/fmsub_b7-01", "37f0",
    "rv32i_m/F/fmsub_b8-01", "13f30",
    "rv32i_m/F/fmul_b1-01", "7220",
    "rv32i_m/F/fmul_b2-01", "38c0",
    "rv32i_m/F/fmul_b3-01", "b320",
    "rv32i_m/F/fmul_b4-01", "3480",
    "rv32i_m/F/fmul_b5-01", "3700",
    "rv32i_m/F/fmul_b6-01", "3480", 
    "rv32i_m/F/fmul_b7-01", "3520",
    "rv32i_m/F/fmul_b8-01", "104a0",
    "rv32i_m/F/fmul_b9-01", "d960",
    "rv32i_m/F/fmv.w.x_b25-01", "2090",
    "rv32i_m/F/fmv.w.x_b26-01", "2090",
    "rv32i_m/F/fmv.x.w_b1-01", "2090",
    "rv32i_m/F/fmv.x.w_b22-01", "2090",
    "rv32i_m/F/fmv.x.w_b23-01", "2090",
    "rv32i_m/F/fmv.x.w_b24-01", "2090",
    "rv32i_m/F/fmv.x.w_b27-01", "2090",
    "rv32i_m/F/fmv.x.w_b28-01", "2090",
    "rv32i_m/F/fmv.x.w_b29-01", "2090",
    "rv32i_m/F/fnmadd_b1-01", "96870",
    "rv32i_m/F/fnmadd_b14-01", "23d0",
// timeconsuming    "rv32i_m/F/fnmadd_b15-01", "19bb40",
    "rv32i_m/F/fnmadd_b16-01", "39d0",
    "rv32i_m/F/fnmadd_b17-01", "39d0",
    "rv32i_m/F/fnmadd_b18-01", "4d10", 
    "rv32i_m/F/fnmadd_b2-01", "4d60",
    "rv32i_m/F/fnmadd_b3-01", "d4f0",
    "rv32i_m/F/fnmadd_b4-01", "3700",
    "rv32i_m/F/fnmadd_b5-01", "3ac0",
    "rv32i_m/F/fnmadd_b6-01", "3700",
    "rv32i_m/F/fnmadd_b7-01", "37f0",
    "rv32i_m/F/fnmadd_b8-01", "13f30",
    "rv32i_m/F/fnmsub_b1-01", "96870",
    "rv32i_m/F/fnmsub_b14-01", "23d0", 
// timeconsuming    "rv32i_m/F/fnmsub_b15-01", "19bb30",
    "rv32i_m/F/fnmsub_b16-01", "39d0",
    "rv32i_m/F/fnmsub_b17-01", "39d0",
    "rv32i_m/F/fnmsub_b18-01", "4d10", 
    "rv32i_m/F/fnmsub_b2-01", "4d60",
    "rv32i_m/F/fnmsub_b3-01", "d4f0",
    "rv32i_m/F/fnmsub_b4-01", "3700",
    "rv32i_m/F/fnmsub_b5-01", "3ac0",
    "rv32i_m/F/fnmsub_b6-01", "3700",
    "rv32i_m/F/fnmsub_b7-01", "37f0", 
    "rv32i_m/F/fnmsub_b8-01", "13f30",
    "rv32i_m/F/fsgnj_b1-01", "7220",
    "rv32i_m/F/fsgnjn_b1-01", "7220",
    "rv32i_m/F/fsgnjx_b1-01", "7220",
    // "rv32i_m/F/fsqrt_b1-01", "2090", // flag i am skiping sqrt
    // "rv32i_m/F/fsqrt_b2-01", "2090",
    // "rv32i_m/F/fsqrt_b20-01", "2090",
    // "rv32i_m/F/fsqrt_b3-01", "2090",
    // "rv32i_m/F/fsqrt_b4-01", "2090",
    // "rv32i_m/F/fsqrt_b5-01", "2090",
    // "rv32i_m/F/fsqrt_b7-01", "2090",
    // "rv32i_m/F/fsqrt_b8-01", "2090",
    // "rv32i_m/F/fsqrt_b9-01", "3310",
    "rv32i_m/F/fsub_b1-01", "7220",
    "rv32i_m/F/fsub_b10-01", "2250",
    "rv32i_m/F/fsub_b11-01", "3fb40",
    "rv32i_m/F/fsub_b12-01", "21b0",
    "rv32i_m/F/fsub_b13-01", "3660",
    "rv32i_m/F/fsub_b2-01", "38b0",
    "rv32i_m/F/fsub_b3-01", "b320",
    "rv32i_m/F/fsub_b4-01", "3480",
    "rv32i_m/F/fsub_b5-01", "3700",
    "rv32i_m/F/fsub_b7-01", "3520", 
    "rv32i_m/F/fsub_b8-01", "104a0",
    "rv32i_m/F/fsw-align-01", "2010"
};


  string arch32c[] = '{
    `RISCVARCHTEST,
    "rv32i_m/C/cadd-01", "4010",
    "rv32i_m/C/caddi-01", "3010",
    "rv32i_m/C/caddi16sp-01", "2010",
    "rv32i_m/C/caddi4spn-01", "2010",
    "rv32i_m/C/cand-01", "4010",
    "rv32i_m/C/candi-01", "3010",
    "rv32i_m/C/cbeqz-01", "3010",
    "rv32i_m/C/cbnez-01", "3010",
    "rv32i_m/C/cj-01", "3010",
    "rv32i_m/C/cjal-01", "3010",
    "rv32i_m/C/cjalr-01", "2010",
    "rv32i_m/C/cjr-01", "2010",
    "rv32i_m/C/cli-01", "2010",
    "rv32i_m/C/clui-01", "2010",
    "rv32i_m/C/clw-01", "2010",
    "rv32i_m/C/clwsp-01", "2010",
    "rv32i_m/C/cmv-01", "2010",
    "rv32i_m/C/cnop-01", "2010",
    "rv32i_m/C/cor-01", "4010",
    "rv32i_m/C/cslli-01", "2010",
    "rv32i_m/C/csrai-01", "2010",
    "rv32i_m/C/csrli-01", "2010",
    "rv32i_m/C/csub-01", "4010",
    "rv32i_m/C/csw-01", "2010",
    "rv32i_m/C/cswsp-01", "2010",
    "rv32i_m/C/cxor-01", "4010"
  };

  string arch32cpriv[] = '{
  //  `RISCVARCHTEST,
      "rv32i_m/C/cebreak-01", "2050"
  };      


  string arch32i[] = '{
    `RISCVARCHTEST,
    "rv32i_m/I/add-01", "5010",
    "rv32i_m/I/addi-01", "4010",
    "rv32i_m/I/and-01", "5010",
    "rv32i_m/I/andi-01", "4010",
    "rv32i_m/I/auipc-01", "2010",
    "rv32i_m/I/beq-01", "39010",
    "rv32i_m/I/bge-01", "3a010",
    "rv32i_m/I/bgeu-01", "4a010",
    "rv32i_m/I/blt-01", "38010",
    "rv32i_m/I/bltu-01", "4b010",
    "rv32i_m/I/bne-01", "39010",
    "rv32i_m/I/fence-01", "2010",
    "rv32i_m/I/jal-01", "1ad010",
    "rv32i_m/I/jalr-01", "2010",
    "rv32i_m/I/lb-align-01", "2010",
    "rv32i_m/I/lbu-align-01", "2010",
    "rv32i_m/I/lh-align-01", "2010",
    "rv32i_m/I/lhu-align-01", "2010",
    "rv32i_m/I/lui-01", "2010",
    "rv32i_m/I/lw-align-01", "2010",
    "rv32i_m/I/or-01", "5010",
    "rv32i_m/I/ori-01", "4010",
    "rv32i_m/I/sb-align-01", "2010",
    "rv32i_m/I/sh-align-01", "2010",
    "rv32i_m/I/sll-01", "2010",
    "rv32i_m/I/slli-01", "2010",
    "rv32i_m/I/slt-01", "5010",
    "rv32i_m/I/slti-01", "4010",
    "rv32i_m/I/sltiu-01", "4010",
    "rv32i_m/I/sltu-01", "5010",
    "rv32i_m/I/sra-01", "2010",
    "rv32i_m/I/srai-01", "2010",
    "rv32i_m/I/srl-01", "2010",
    "rv32i_m/I/srli-01", "2010",
    "rv32i_m/I/sub-01", "5010",
    "rv32i_m/I/sw-align-01", "2010",
    "rv32i_m/I/xor-01", "5010",
    "rv32i_m/I/xori-01", "4010"
  };

 string wally64i[] = '{
    `WALLYTEST,
    "rv64i_m/I/WALLY-ADD", "002010",
    "rv64i_m/I/WALLY-SLT", "002010",
    "rv64i_m/I/WALLY-SLTU", "002010",
    "rv64i_m/I/WALLY-SUB", "002010",
    "rv64i_m/I/WALLY-XOR", "002010"
 };

 string wally64priv[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-CSR-permission-s-01", "0060a0",
    //"rv64i_m/privilege/WALLY-CSR-PERMISSIONS-M", "005090",
    //"rv64i_m/privilege/WALLY-CSR-PERMISSIONS-S", "003090",
    "rv64i_m/privilege/WALLY-CSR-permission-u-01", "0060a0",
   // "rv64i_m/privilege/WALLY-MARCHID", "004090",
/*    "rv64i_m/privilege/WALLY-MCAUSE", "003090",
    "rv64i_m/privilege/WALLY-MEDELEG", "004090",
    "rv64i_m/privilege/WALLY-MHARTID", "004090",
    "rv64i_m/privilege/WALLY-MIMPID", "004090",*/
    "rv64i_m/privilege/WALLY-minfo-01", "0050a0",
    "rv64i_m/privilege/WALLY-misa-01", "0050a0",
    "rv64i_m/privilege/WALLY-MMU-SV39", "0050a0",
    "rv64i_m/privilege/WALLY-MMU-SV48", "0050a0",
/*    "rv64i_m/privilege/WALLY-MSTATUS", "002090",
    "rv64i_m/privilege/WALLY-MTVEC", "002090",
    "rv64i_m/privilege/WALLY-MVENDORID", "004090", */
    "rv64i_m/privilege/WALLY-PMA", "0050a0",
    "rv64i_m/privilege/WALLY-PMP", "0050a0",
//    "rv64i_m/privilege/WALLY-SCAUSE", "002090",
//    "rv64i_m/privilege/WALLY-scratch-01", "0040a0",
//    "rv64i_m/privilege/WALLY-sscratch-s-01", "0040a0",
    "rv64i_m/privilege/WALLY-trap-01", "0050a0",
    "rv64i_m/privilege/WALLY-trap-s-01", "0050a0",
    "rv64i_m/privilege/WALLY-trap-u-01", "0050a0",
    "rv64i_m/privilege/WALLY-MIE-01", "0050a0",
    "rv64i_m/privilege/WALLY-mtvec-01", "0050a0",
    "rv64i_m/privilege/WALLY-stvec-01", "0050a0",
    "rv64i_m/privilege/WALLY-PIE-stack-01", "0050a0",
    "rv64i_m/privilege/WALLY-PIE-stack-s-01", "0050a0",
    "rv64i_m/privilege/WALLY-trap-sret-01", "0050a0"
    // "rv64i_m/privilege/WALLY-status-tw-01", "0050a0",
    // "rv64i_m/privilege/WALLY-WFI-01", "0050a0",
    // "rv64i_m/privilege/WALLY-status-fp-01", "0050a0"
//    "rv64i_m/privilege/WALLY-STVEC", "002090",
//    "rv64i_m/privilege/WALLY-UCAUSE", "002090",

 };

 string wally64periph[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-PERIPH", "3310"
 };

 string wally32e[] = '{
    `WALLYTEST,
    "rv32i_m/I/E-beq-01", "03b010",
    "rv32i_m/I/E-add-01", "005010",
    "rv32i_m/I/E-addi-01", "004010",
    "rv32i_m/I/E-and-01", "005010",
    "rv32i_m/I/E-andi-01", "004010",
    "rv32i_m/I/E-auipc-01", "002010",
    "rv32i_m/I/E-bge-01", "034010",
    "rv32i_m/I/E-bgeu-01", "047010",
    "rv32i_m/I/E-blt-01", "038010",
    "rv32i_m/I/E-bltu-01", "03e010",
    "rv32i_m/I/E-bne-01", "038010",
    "rv32i_m/I/E-jal-01", "e02010",
    "rv32i_m/I/E-jalr-01", "002010",
    "rv32i_m/I/E-lb-align-01", "002010",
    "rv32i_m/I/E-lbu-align-01", "002010",
    "rv32i_m/I/E-lh-align-01", "002010",
    "rv32i_m/I/E-lhu-align-01", "002010",
    "rv32i_m/I/E-lui-01", "002010",
    "rv32i_m/I/E-lw-align-01", "002010",
    "rv32i_m/I/E-or-01", "005010",
    "rv32i_m/I/E-ori-01", "004010",
    "rv32i_m/I/E-sb-align-01", "002010",
    "rv32i_m/I/E-sh-align-01", "002010",
    "rv32i_m/I/E-sll-01", "002010",
    "rv32i_m/I/E-slli-01", "002010",
    "rv32i_m/I/E-slt-01", "005010",
    "rv32i_m/I/E-slti-01", "004010",
    "rv32i_m/I/E-sltiu-01", "004010",
    "rv32i_m/I/E-sltu-01", "005010",
    "rv32i_m/I/E-sra-01", "002010",
    "rv32i_m/I/E-srai-01", "002010",
    "rv32i_m/I/E-srl-01", "002010",
    "rv32i_m/I/E-srli-01", "002010",
    "rv32i_m/I/E-sub-01", "005010",
    "rv32i_m/I/E-sw-align-01", "002010",
    "rv32i_m/I/E-xor-01", "005010",
    "rv32i_m/I/E-xori-01", "004010"
 };

string wally32i[] = '{
    `WALLYTEST,
    "rv32i_m/I/WALLY-ADD", "002010",
    "rv32i_m/I/WALLY-SLT", "002010",
    "rv32i_m/I/WALLY-SLTU", "002010",
    "rv32i_m/I/WALLY-SUB", "002010",
    "rv32i_m/I/WALLY-XOR", "002010"
 };

 string wally32priv[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/WALLY-CSR-permission-s-01", "006080",
    "rv32i_m/privilege/WALLY-CSR-permission-u-01", "006080",
    "rv32i_m/privilege/WALLY-minfo-01", "005080",
    "rv32i_m/privilege/WALLY-misa-01", "005080",
    "rv32i_m/privilege/WALLY-MMU-SV32", "005080",
    "rv32i_m/privilege/WALLY-PMA", "005080",
    "rv32i_m/privilege/WALLY-PMP", "005080",
    "rv32i_m/privilege/WALLY-trap-01", "005080",
    "rv32i_m/privilege/WALLY-trap-s-01", "005080",
    "rv32i_m/privilege/WALLY-trap-u-01", "005080",
    "rv32i_m/privilege/WALLY-MIE-01", "005080",
    "rv32i_m/privilege/WALLY-mtvec-01", "005080",
    "rv32i_m/privilege/WALLY-stvec-01", "005080",
    "rv32i_m/privilege/WALLY-PIE-stack-01", "005080",
    "rv32i_m/privilege/WALLY-PIE-stack-s-01", "005080",
    "rv32i_m/privilege/WALLY-trap-sret-01", "005080"

 };

 string wally32periph[] = '{
    `WALLYTEST
 };



// Populate parameter structure with values specific to the current configuration

parameter cvw_t P = '{ 
  FPGA :        FPGA,  
  QEMU :         QEMU,  
  XLEN :         XLEN,  
  IEEE754 :        IEEE754, 
  MISA : MISA, 
  AHBW :         AHBW, 
  ZICSR_SUPPORTED :        ZICSR_SUPPORTED,
  ZIFENCEI_SUPPORTED :        ZIFENCEI_SUPPORTED,
  COUNTERS :         COUNTERS,
  ZICOUNTERS_SUPPORTED :        ZICOUNTERS_SUPPORTED,
  ZFH_SUPPORTED :        ZFH_SUPPORTED,
  SSTC_SUPPORTED :        SSTC_SUPPORTED,
  VIRTMEM_SUPPORTED :        VIRTMEM_SUPPORTED,
  VECTORED_INTERRUPTS_SUPPORTED :        VECTORED_INTERRUPTS_SUPPORTED,
  BIGENDIAN_SUPPORTED :        BIGENDIAN_SUPPORTED,
  SVADU_SUPPORTED :        SVADU_SUPPORTED,
  ZMMUL_SUPPORTED :        ZMMUL_SUPPORTED,
  BUS_SUPPORTED :        BUS_SUPPORTED,
  DCACHE_SUPPORTED :        DCACHE_SUPPORTED,
  ICACHE_SUPPORTED :        ICACHE_SUPPORTED,
  ITLB_ENTRIES :        ITLB_ENTRIES,
  DTLB_ENTRIES :        DTLB_ENTRIES,
  DCACHE_NUMWAYS :        DCACHE_NUMWAYS,
  DCACHE_WAYSIZEINBYTES :        DCACHE_WAYSIZEINBYTES,
  DCACHE_LINELENINBITS :        DCACHE_LINELENINBITS,
  ICACHE_NUMWAYS :        ICACHE_NUMWAYS,
  ICACHE_WAYSIZEINBYTES :        ICACHE_WAYSIZEINBYTES,
  ICACHE_LINELENINBITS :        ICACHE_LINELENINBITS,
  IDIV_BITSPERCYCLE :        IDIV_BITSPERCYCLE,
  IDIV_ON_FPU :        IDIV_ON_FPU,
  PMP_ENTRIES :        PMP_ENTRIES,
  RESET_VECTOR :        RESET_VECTOR,
  WFI_TIMEOUT_BIT :        WFI_TIMEOUT_BIT,
  DTIM_SUPPORTED :        DTIM_SUPPORTED,
  DTIM_BASE :        DTIM_BASE,
  DTIM_RANGE :        DTIM_RANGE,
  IROM_SUPPORTED :        IROM_SUPPORTED,
  IROM_BASE :        IROM_BASE,
  IROM_RANGE :        IROM_RANGE,
  BOOTROM_SUPPORTED :        BOOTROM_SUPPORTED,
  BOOTROM_BASE :        BOOTROM_BASE,
  BOOTROM_RANGE :        BOOTROM_RANGE,
  UNCORE_RAM_SUPPORTED :        UNCORE_RAM_SUPPORTED,
  UNCORE_RAM_BASE :        UNCORE_RAM_BASE,
  UNCORE_RAM_RANGE :        UNCORE_RAM_RANGE,
  EXT_MEM_SUPPORTED :        EXT_MEM_SUPPORTED,
  EXT_MEM_BASE :        EXT_MEM_BASE,
  EXT_MEM_RANGE :        EXT_MEM_RANGE,
  CLINT_SUPPORTED :        CLINT_SUPPORTED,
  CLINT_BASE :        CLINT_BASE,
  CLINT_RANGE :        CLINT_RANGE,
  GPIO_SUPPORTED :        GPIO_SUPPORTED,
  GPIO_BASE :        GPIO_BASE,
  GPIO_RANGE :        GPIO_RANGE,
  UART_SUPPORTED :        UART_SUPPORTED,
  UART_BASE :        UART_BASE,
  UART_RANGE :        UART_RANGE,
  PLIC_SUPPORTED :        PLIC_SUPPORTED,
  PLIC_BASE :        PLIC_BASE,
  PLIC_RANGE :        PLIC_RANGE,
  SDC_SUPPORTED :        SDC_SUPPORTED,
  SDC_BASE :        SDC_BASE,
  SDC_RANGE :        SDC_RANGE,
  GPIO_LOOPBACK_TEST :        GPIO_LOOPBACK_TEST,
  UART_PRESCALE :        UART_PRESCALE ,
  PLIC_NUM_SRC :        PLIC_NUM_SRC,
  PLIC_NUM_SRC_LT_32 :        PLIC_NUM_SRC_LT_32,
  PLIC_GPIO_ID :        PLIC_GPIO_ID,
  PLIC_UART_ID :        PLIC_UART_ID,
  BPRED_SUPPORTED :        BPRED_SUPPORTED,
  //parameter :        BPRED_TYPE "BP_GSHARE" // BP_GSHARE_BASIC, BP_GLOBAL, BP_GLOBAL_BASIC, BP_TWOBIT
  BPRED_SIZE :        BPRED_SIZE,
  BTB_SIZE :        BTB_SIZE,
  RADIX :        RADIX,
  DIVCOPIES :        DIVCOPIES,
  ZBA_SUPPORTED :        ZBA_SUPPORTED,
  ZBB_SUPPORTED :        ZBB_SUPPORTED,
  ZBC_SUPPORTED :        ZBC_SUPPORTED,
  ZBS_SUPPORTED :        ZBS_SUPPORTED,
  A_SUPPORTED :        A_SUPPORTED,
  B_SUPPORTED :        B_SUPPORTED,
  C_SUPPORTED :        C_SUPPORTED,
  D_SUPPORTED :        D_SUPPORTED,
  E_SUPPORTED :        E_SUPPORTED,
  F_SUPPORTED :        F_SUPPORTED,
  I_SUPPORTED :        I_SUPPORTED,
  M_SUPPORTED :        M_SUPPORTED,
  Q_SUPPORTED :        Q_SUPPORTED,
  S_SUPPORTED :        S_SUPPORTED,
  U_SUPPORTED :        U_SUPPORTED,
  USE_SRAM :        USE_SRAM,
  LLEN :LLEN,
  FLEN :FLEN,
  VPN_SEGMENT_BITS :VPN_SEGMENT_BITS,
  PA_BITS :         PA_BITS
};

///////////////////////////////////////////
// irom.sv
//
// Written: Ross Thompson ross1728@gmail.com January 30, 2022
// Modified: 
//
// Purpose: simple instruction ROM
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// MIT LICENSE
// Permission is hereby granted, free of charge, to any person obtaining a copy of this 
// software and associated documentation files (the "Software"), to deal in the Software 
// without restriction, including without limitation the rights to use, copy, modify, merge, 
// publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons 
// to whom the Software is furnished to do so, subject to the following conditions:
//
//   The above copyright notice and this permission notice shall be included in all copies or 
//   substantial portions of the Software.
//
//   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, 
//   INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR 
//   PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS 
//   BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, 
//   TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE 
//   OR OTHER DEALINGS IN THE SOFTWARE.
////////////////////////////////////////////////////////////////////////////////////////////////

`include "wally-config.vh"

module irom(
  input logic               clk, reset, ce,
  input logic [`XLEN-1:0]   Adr,
  output logic [31:0]  ReadData
);

  localparam ADDR_WDITH = $clog2(`IROM_RANGE/8); 
  localparam OFFSET = $clog2(`XLEN/8);

  logic [`XLEN-1:0] ReadDataFull;

  rom1p1r #(ADDR_WDITH, `XLEN) rom(.clk, .ce, .addr(Adr[ADDR_WDITH+OFFSET-1:OFFSET]), .dout(ReadDataFull));
  if (`XLEN == 32) begin
	logic AdrD;
    flopen #(1) AdrReg(clk, ce, Adr[1], AdrD);
	assign ReadData = AdrD ? {16'b0, ReadDataFull[31:16]} : ReadDataFull;
  end
  // have to delay Ardr[OFFSET-1] by 1 cycle
  else             begin
    logic [OFFSET-2:0] AdrD;
    flopen #(OFFSET-1) AdrReg(clk, ce, Adr[OFFSET-1:1], AdrD);
    assign ReadData = AdrD == 2'b11 ? {16'b0, ReadDataFull[63:48]} :
					  AdrD == 2'b10 ? ReadDataFull[63:32] :
					  AdrD == 2'b01 ? ReadDataFull[47:16] :
					  ReadDataFull[31:0];
  end
endmodule  
  

///////////////////////////////////////////
// tests.vh
//
// Written: David_Harris@hmc.edu 7 October 2021
// Modified:
//
// Purpose: List of tests to apply
//
// A component of the Wally configurable RISC-V project.
//
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define RISCVARCHTEST "0"
`define WALLYTEST "1"
`define COREMARK "2"
`define EMBENCH "3"
`define CUSTOM "4"
`define COVERAGE "5"
`define BUILDROOT "6"

string tvpaths[] = '{
  "../../tests/riscof/work/riscv-arch-test/",
  "../../tests/riscof/work/wally-riscv-arch-test/",
  "../../benchmarks/coremark/work/",
  "../../addins/embench-iot/",
  "../../tests/custom/work/",
  "../../tests/coverage/"
};

string coverage64gc[] = '{
  `COVERAGE,
  "ieu",
  "priv",
  "ebu",
  "csrwrites",
  "ifu",
  "fpu",
  "lsu",
  "vm64check",
  "tlbmisc",
  "tlbNAPOT",
  "tlbASID",
  "tlbGLB",
  "tlbMP",
  "tlbGP",
  "tlbTP",
  "tlbMisaligned",
  "hptwAccessFault",
  "nonleafpbmtfault",
  "amoAccessFault",
  "floatmisc",
  "ifuCamlineWrite",
  "dcache1",
  "dcache2",
  "pmp",
  "pmpcfg",
  "pmpcfg1",
  "pmpcfg2",
  "pmppriority",
  "pmpcbo",
  "pmpadrdecs",
  "btbthrash"
};

string buildroot[] = '{
  `BUILDROOT,
  "buildroot"
};

string coremark[] = '{
  `COREMARK,
  "coremark.bare.riscv"
};

string embench[] = '{
  `EMBENCH,
  "bd_speedopt_speed/src/aha-mont64/aha-mont64",
  "bd_speedopt_speed/src/crc32/crc32",
  "bd_speedopt_speed/src/cubic/cubic", // cubic is likely going to removed when embench 2.0 launches
  "bd_speedopt_speed/src/edn/edn",
  "bd_speedopt_speed/src/huffbench/huffbench",
  "bd_speedopt_speed/src/matmult-int/matmult-int",
  "bd_speedopt_speed/src/md5sum/md5sum", //commenting out tests from embench 2.0. When embench 2.0 launches stably, add these tests back
  "bd_speedopt_speed/src/minver/minver",
  "bd_speedopt_speed/src/nettle-aes/nettle-aes",
  "bd_speedopt_speed/src/nettle-sha256/nettle-sha256",
  "bd_speedopt_speed/src/nsichneu/nsichneu",
  "bd_speedopt_speed/src/nbody/nbody",
  "bd_speedopt_speed/src/picojpeg/picojpeg",
  "bd_speedopt_speed/src/primecount/primecount",
  "bd_speedopt_speed/src/qrduino/qrduino",
  "bd_speedopt_speed/src/sglib-combined/sglib-combined",
  "bd_speedopt_speed/src/slre/slre",
  "bd_speedopt_speed/src/st/st",
  "bd_speedopt_speed/src/statemate/statemate",
  "bd_speedopt_speed/src/tarfind/tarfind",
  "bd_speedopt_speed/src/ud/ud",
  "bd_speedopt_speed/src/wikisort/wikisort",
  "bd_sizeopt_speed/src/aha-mont64/aha-mont64",
  "bd_sizeopt_speed/src/crc32/crc32",
  "bd_sizeopt_speed/src/cubic/cubic",
  "bd_sizeopt_speed/src/edn/edn",
  "bd_sizeopt_speed/src/huffbench/huffbench",
  "bd_sizeopt_speed/src/matmult-int/matmult-int",
  "bd_sizeopt_speed/src/md5sum/md5sum",
  "bd_sizeopt_speed/src/minver/minver",
  "bd_sizeopt_speed/src/nbody/nbody",
  "bd_sizeopt_speed/src/nettle-aes/nettle-aes",
  "bd_sizeopt_speed/src/nettle-sha256/nettle-sha256",
  "bd_sizeopt_speed/src/nsichneu/nsichneu",
  "bd_sizeopt_speed/src/picojpeg/picojpeg",
  "bd_sizeopt_speed/src/primecount/primecount",
  "bd_sizeopt_speed/src/qrduino/qrduino",
  "bd_sizeopt_speed/src/sglib-combined/sglib-combined",
  "bd_sizeopt_speed/src/slre/slre",
  "bd_sizeopt_speed/src/st/st",
  "bd_sizeopt_speed/src/statemate/statemate",
  "bd_sizeopt_speed/src/tarfind/tarfind",
  "bd_sizeopt_speed/src/ud/ud",
  "bd_sizeopt_speed/src/wikisort/wikisort"
};

string wally64q[] = '{
  `WALLYTEST,
  "rv64i_m/Q/src/WALLY-q-01.S"
};

string wally64a_lrsc[] = '{
  `WALLYTEST,
  "rv64i_m/privilege/src/WALLY-lrsc-01.S"
};

string wally32a_lrsc[] = '{
  `WALLYTEST,
  "rv32i_m/privilege/src/WALLY-lrsc-01.S"
};

string arch32pmp[] = '{
  `RISCVARCHTEST,
  "rv32i_m/pmp/src/pmpf_cfg_wr.S",
  "rv32i_m/pmp/src/pmpm_cfg_A_all.S",
  "rv32i_m/pmp/src/pmpm_cfg_A_off_all.S",
  "rv32i_m/pmp/src/pmpm_cfg_A_tor_bot.S",
  "rv32i_m/pmp/src/pmpm_cfg_A_tor_zero.S",
  "rv32i_m/pmp/src/pmpm_cfg_L_access_all.S",
  "rv32i_m/pmp/src/pmpm_cfg_L_modify_napot.S",
  "rv32i_m/pmp/src/pmpm_cfg_L_modify_off.S",
  "rv32i_m/pmp/src/pmpm_cfg_L_modify_tor.S",
  "rv32i_m/pmp/src/pmpm_cfg_XWR_all-01.S",
  "rv32i_m/pmp/src/pmpm_cfg_XWR_all-02.S",
  "rv32i_m/pmp/src/pmpm_cfg_XWR_all-03.S",
  "rv32i_m/pmp/src/pmpm_cfg_XWR_all-04.S",
  "rv32i_m/pmp/src/pmpm_cfg_napot_all.S",
  "rv32i_m/pmp/src/pmpm_cfg_tor_all.S",
  "rv32i_m/pmp/src/pmpm_cfg_tor_check-01.S",
  "rv32i_m/pmp/src/pmpm_cfg_tor_check-02.S",
  "rv32i_m/pmp/src/pmpm_cfg_tor_check-03.S",
  "rv32i_m/pmp/src/pmpm_grain.S",
  "rv32i_m/pmp/src/pmpm_grain_check.S",
  "rv32i_m/pmp/src/pmpm_misaligned_napot.S",
  "rv32i_m/pmp/src/pmpm_misaligned_off.S",
  "rv32i_m/pmp/src/pmpm_misaligned_tor.S",
  "rv32i_m/pmp/src/pmpm_napot_legal_lwxr.S",
  "rv32i_m/pmp/src/pmpm_priority.S",
  "rv32i_m/pmp/src/pmpm_priority_off.S",
  "rv32i_m/pmp/src/pmpm_tor_legal_lwxr.S",
  "rv32i_m/pmp/src/pmps_cfg_A_off.S",
  "rv32i_m/pmp/src/pmps_cfg_XWR.S",
  "rv32i_m/pmp/src/pmps_csr_access.S",
  "rv32i_m/pmp/src/pmps_mprv_check-01.S",
  "rv32i_m/pmp/src/pmps_mprv_check-02.S",
  "rv32i_m/pmp/src/pmps_napot_legal_lxwr.S",
  "rv32i_m/pmp/src/pmps_none.S",
  "rv32i_m/pmp/src/pmps_tor_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpu_cfg_A_off.S",
  "rv32i_m/pmp/src/pmpu_cfg_XWR.S",
  "rv32i_m/pmp/src/pmpu_csr_access.S",
  "rv32i_m/pmp/src/pmpu_mprv_check-01.S",
  "rv32i_m/pmp/src/pmpu_mprv_check-02.S",
  "rv32i_m/pmp/src/pmpu_napot_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpu_none.S",
  "rv32i_m/pmp/src/pmpu_tor_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpzaamo_cfg_wr.S",
  "rv32i_m/pmp/src/pmpzca_aligned_napot.S",
  "rv32i_m/pmp/src/pmpzca_aligned_off.S",
  "rv32i_m/pmp/src/pmpzca_aligned_tor.S",
  "rv32i_m/pmp/src/pmpzca_cret_napot.S",
  "rv32i_m/pmp/src/pmpzca_cret_tor.S",
  "rv32i_m/pmp/src/pmpzca_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpzca_misaligned_napot.S",
  "rv32i_m/pmp/src/pmpzca_misaligned_off.S",
  "rv32i_m/pmp/src/pmpzca_misaligned_tor.S",
  "rv32i_m/pmp/src/pmpzcb_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpzcd_legal_lxwr.S",
  "rv32i_m/pmp/src/pmpzcf_legal_lxwr.S"
  // *** Uncomment following when G = 0
  //"rv32i_m/pmp/src/pmpzca_misaligned_na4.S",
  //"rv32i_m/pmp/src/pmpzca_cret_na4.S",
  //"rv32i_m/pmp/src/pmpzca_aligned_na4.S",
  //"rv32i_m/pmp/src/pmpu_na4_legal_lxwr.S",
  //"rv32i_m/pmp/src/pmps_na4_legal_lxwr.S",
  //"rv32i_m/pmp/src/pmpm_na4_legal_lwxr.S",
  //"rv32i_m/pmp/src/pmpm_misaligned_na4.S",
  //"rv32i_m/pmp/src/pmpm_cfg_na4_all.S",
  // *** Uncomment following when PMP Entries = 64
  //"rv32i_m/pmp/src/pmpm_all_entries_check-01.S",  
  //"rv32i_m/pmp/src/pmpm_all_entries_check-02.S",
  //"rv32i_m/pmp/src/pmpm_all_entries_check-03.S",
  //"rv32i_m/pmp/src/pmpm_all_entries_check-04.S",
  // *** Uncomment following when PR#705 is merged
  //"rv32i_m/pmp/src/pmpm_csr_walk.S",
  //"rv32i_m/pmp/src/pmpzicbo_prefetch.S",
  // *** Uncomment following when PR#699 is merged
  //"rv32i_m/pmp/src/pmpzicbo_cbo_WR_01.S",  
  //"rv32i_m/pmp/src/pmpzicbo_cbo_WR_02.S",
  //"rv32i_m/pmp/src/pmpzicbo_cbo_WR_03.S",
  //"rv32i_m/pmp/src/pmpzalrsc_cfg_wr.S"
};

string arch64pmp[] = '{
  `RISCVARCHTEST,
  "rv64i_m/pmp/src/pmpf_cfg_wr.S",
  "rv64i_m/pmp/src/pmpm_cfg_A_all.S",
  "rv64i_m/pmp/src/pmpm_cfg_A_off_all.S",
  "rv64i_m/pmp/src/pmpm_cfg_A_tor_bot.S",
  "rv64i_m/pmp/src/pmpm_cfg_A_tor_zero.S",
  "rv64i_m/pmp/src/pmpm_cfg_L_access_all.S",
  "rv64i_m/pmp/src/pmpm_cfg_L_modify_napot.S",
  "rv64i_m/pmp/src/pmpm_cfg_L_modify_off.S",
  "rv64i_m/pmp/src/pmpm_cfg_L_modify_tor.S",
  "rv64i_m/pmp/src/pmpm_cfg_XWR_all-01.S",
  "rv64i_m/pmp/src/pmpm_cfg_XWR_all-02.S",
  "rv64i_m/pmp/src/pmpm_cfg_XWR_all-03.S",
  "rv64i_m/pmp/src/pmpm_cfg_XWR_all-04.S",
  "rv64i_m/pmp/src/pmpm_cfg_napot_all.S",
  "rv64i_m/pmp/src/pmpm_cfg_tor_all.S",
  "rv64i_m/pmp/src/pmpm_cfg_tor_check-01.S",
  "rv64i_m/pmp/src/pmpm_cfg_tor_check-02.S",
  "rv64i_m/pmp/src/pmpm_cfg_tor_check-03.S",
  "rv64i_m/pmp/src/pmpm_csr_walk.S",
  "rv64i_m/pmp/src/pmpm_grain.S",
  "rv64i_m/pmp/src/pmpm_grain_check.S",
  "rv64i_m/pmp/src/pmpm_napot_legal_lxwr.S",
  "rv64i_m/pmp/src/pmpm_priority.S",
  "rv64i_m/pmp/src/pmpm_priority_off.S",
  "rv64i_m/pmp/src/pmpm_tor_legal_lxwr.S",
  "rv64i_m/pmp/src/pmps_cfg_A_off.S",
  "rv64i_m/pmp/src/pmps_cfg_XWR.S",
  "rv64i_m/pmp/src/pmps_csr_access.S",
  "rv64i_m/pmp/src/pmps_mprv_check-01.S",
  "rv64i_m/pmp/src/pmps_mprv_check-02.S",
  "rv64i_m/pmp/src/pmps_napot_legal_lxwr.S",
  "rv64i_m/pmp/src/pmps_none.S",
  "rv64i_m/pmp/src/pmps_tor_legal_lxwr.S",
  "rv64i_m/pmp/src/pmpu_cfg_A_off.S",
  "rv64i_m/pmp/src/pmpu_cfg_XWR.S",
  "rv64i_m/pmp/src/pmpu_csr_access.S",
  "rv64i_m/pmp/src/pmpu_mprv_check-01.S",
  "rv64i_m/pmp/src/pmpu_mprv_check-02.S",
  "rv64i_m/pmp/src/pmpu_napot_legal_lxwr.S",
  "rv64i_m/pmp/src/pmpu_none.S",
  "rv64i_m/pmp/src/pmpu_tor_legal_lxwr.S",
  "rv64i_m/pmp/src/pmpzaamo_cfg_wr.S",
  "rv64i_m/pmp/src/pmpzca_aligned_napot.S",
  "rv64i_m/pmp/src/pmpzca_aligned_off.S",
  "rv64i_m/pmp/src/pmpzca_aligned_tor.S",
  "rv64i_m/pmp/src/pmpzca_cret_napot.S",
  "rv64i_m/pmp/src/pmpzca_cret_tor.S",
  "rv64i_m/pmp/src/pmpzca_legal_lwxr.S",
  "rv64i_m/pmp/src/pmpzca_misaligned_napot.S",
  "rv64i_m/pmp/src/pmpzca_misaligned_off.S",
  "rv64i_m/pmp/src/pmpzca_misaligned_tor.S",
  "rv64i_m/pmp/src/pmpzcb_legal_lwxr.S",
  "rv64i_m/pmp/src/pmpzcd_legal_lwxr.S"
  // *** Uncomment following when PMP Entries = 64
  //"rv64i_m/pmp/src/pmpm_all_entries_check-01.S",  
  //"rv64i_m/pmp/src/pmpm_all_entries_check-02.S",
  //"rv64i_m/pmp/src/pmpm_all_entries_check-03.S",
  //"rv64i_m/pmp/src/pmpm_all_entries_check-04.S",
  // *** Uncomment following when G = 0
  //"rv64i_m/pmp/src/pmpm_access_double_region.S",
  //"rv64i_m/pmp/src/pmpm_cfg_na4_all.S",
  //"rv64i_m/pmp/src/pmpm_na4_boundary-01.S",
  //"rv64i_m/pmp/src/pmpm_na4_boundary-02.S",
  //"rv64i_m/pmp/src/pmpm_na4_legal_lxwr.S",
  //"rv64i_m/pmp/src/pmpm_tor_boundary-01.S",
  //"rv64i_m/pmp/src/pmpm_tor_boundary-02.S",
  //"rv64i_m/pmp/src/pmps_na4_legal_lxwr.S",
  //"rv64i_m/pmp/src/pmpu_na4_legal_lxwr.S",
  //"rv64i_m/pmp/src/pmpzca_aligned_na4.S",
  //"rv64i_m/pmp/src/pmpzca_cret_na4.S",
  //"rv64i_m/pmp/src/pmpzca_misaligned_na4.S",
  // *** Uncomment following when PR#705 is merged
  //"rv64i_m/pmp/src/pmpzicbo_prefetch.S",
  // *** Uncomment following when PR#699 is merged
  //"rv64i_m/pmp/src/pmpzicbo_cbo_WR_01.S",  
  //"rv64i_m/pmp/src/pmpzicbo_cbo_WR_02.S",
  //"rv64i_m/pmp/src/pmpzicbo_cbo_WR_03.S",
  //"rv64i_m/pmp/src/pmpzalrsc_cfg_wr.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_na4.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_napot.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_tor.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_off.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_na4_wrap.S",
  //"rv64i_m/pmp/src/pmpm_misaligned_tor_wrap.S"
};

string arch32vm_sv32[] = '{
  `RISCVARCHTEST,
  "rv32i_m/vm_sv32/src/mstatus_tvm_test.S",
  "rv32i_m/vm_sv32/src/satp_access_tests.S",
  "rv32i_m/vm_sv32/src/vm_A_and_D_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_A_and_D_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_U_Bit_set_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_U_Bit_unset_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_U_Bit_unset_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_VA_all_ones_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_VA_all_zeros_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_global_pte_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_global_pte_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_invalid_pte_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_invalid_pte_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_misaligned_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_misaligned_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_mprv_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_mprv_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_mprv_U_set_sum_set_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_mprv_U_set_sum_unset_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_mprv_bare_mode.S",
  // "rv32i_m/vm_sv32/src/vm_mstatus_sbe_set_S_mode.S", TODO: Reenable when Sail big endian support is merged
  // "rv32i_m/vm_sv32/src/vm_mstatus_sbe_set_sum_set_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_mxr_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_mxr_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_nleaf_pte_level0_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_nleaf_pte_level0_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_reserved_rsw_pte_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_reserved_rsw_pte_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_reserved_rwx_pte_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_reserved_rwx_pte_U_mode.S",
  "rv32i_m/vm_sv32/src/vm_sum_set_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_sum_set_U_Bit_unset_S_mode.S",
  "rv32i_m/vm_sv32/src/vm_sum_unset_S_mode.S",
  "rv32i_m/vm_pmp/src/sv32_pmp_on_pa_S_mode.S",
  "rv32i_m/vm_pmp/src/sv32_pmp_on_pa_U_mode.S",
  "rv32i_m/vm_pmp/src/sv32_pmp_on_pte_S_mode.S",
  "rv32i_m/vm_pmp/src/sv32_pmp_on_pte_U_mode.S"
};

string arch64vm_sv39[] = '{
  `RISCVARCHTEST,
  "rv64i_m/vm_sv39/src/vm_A_and_D_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_A_and_D_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_VA_all_ones_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_VA_all_zeros_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_canonical_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_canonical_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_res_global_pte_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_res_global_pte_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_invalid_pte_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_invalid_pte_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_misaligned_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_misaligned_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_mprv_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_mprv_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_mprv_U_set_sum_set_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_mprv_U_set_sum_unset_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_mprv_bare_mode.S",
  //"rv64i_m/vm_sv39/src/vm_mstatus_sbe_set_S_mode.S",
  //"rv64i_m/vm_sv39/src/vm_mstatus_sbe_set_sum_set_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_mstatus_tvm_test.S",
  "rv64i_m/vm_sv39/src/vm_mxr_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_mxr_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_nleaf_pte_level0_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_nleaf_pte_level0_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_pte_reserved_field_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_reserved_rsw_pte_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_reserved_rsw_pte_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_reserved_rwx_pte_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_reserved_rwx_pte_U_mode.S",
  //"rv64i_m/vm_sv39/src/vm_reserved_svnapot_S_mode.S",  // Run this if SVNAPOT_SUPPORTED == 0
  "rv64i_m/vm_sv39/src/vm_reserved_svpbmt_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_satp_access_tests.S",
  "rv64i_m/vm_sv39/src/vm_spage_access_U_mode.S",
  "rv64i_m/vm_sv39/src/vm_sum_set_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_sum_set_U_bit_unset_S_mode.S",
  "rv64i_m/vm_sv39/src/vm_sum_unset_S_mode.S",
  "rv64i_m/vm_pmp/src/sv39/sv39_pmp_on_pa_S_mode.S",
  "rv64i_m/vm_pmp/src/sv39/sv39_pmp_on_pa_U_mode.S",
  "rv64i_m/vm_pmp/src/sv39/sv39_pmp_on_pte_S_mode.S",
  "rv64i_m/vm_pmp/src/sv39/sv39_pmp_on_pte_U_mode.S"
};

string arch64vm_sv48[] = '{
  `RISCVARCHTEST,
  "rv64i_m/vm_sv48/src/sv48_A_and_D_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_A_and_D_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_VA_all_ones_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_VA_all_zeros_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_canonical_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_canonical_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_res_global_pte_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_res_global_pte_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_invalid_pte_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_invalid_pte_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_misaligned_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_misaligned_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mprv_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mprv_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mprv_U_set_sum_set_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mprv_U_set_sum_unset_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mprv_bare_mode.S",
  //"rv64i_m/vm_sv48/src/sv48_mstatus_sbe_set_S_mode.S",
  //"rv64i_m/vm_sv48/src/sv48_mstatus_sbe_set_sum_set_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mstatus_tvm_test.S",
  "rv64i_m/vm_sv48/src/sv48_mxr_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_mxr_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_nleaf_pte_level0_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_nleaf_pte_level0_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_pte_reserved_field_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_reserved_rsw_pte_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_reserved_rsw_pte_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_reserved_rwx_pte_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_reserved_rwx_pte_U_mode.S",
  //"rv64i_m/vm_sv48/src/sv48_reserved_svnapot_S_mode.S",  // Run this if SVNAPOT_SUPPORTED == 0
  "rv64i_m/vm_sv48/src/sv48_reserved_svpbmt_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_satp_access_tests.S",
  "rv64i_m/vm_sv48/src/sv48_spage_access_U_mode.S",
  "rv64i_m/vm_sv48/src/sv48_sum_set_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_sum_set_U_bit_unset_S_mode.S",
  "rv64i_m/vm_sv48/src/sv48_sum_unset_S_mode.S",
  "rv64i_m/vm_pmp/src/sv48/sv48_pmp_on_pa_S_mode.S",
  "rv64i_m/vm_pmp/src/sv48/sv48_pmp_on_pa_U_mode.S",
  "rv64i_m/vm_pmp/src/sv48/sv48_pmp_on_pte_S_mode.S",
  "rv64i_m/vm_pmp/src/sv48/sv48_pmp_on_pte_U_mode.S"
};

string arch64priv[] = '{
  `RISCVARCHTEST,
  "rv64i_m/privilege/src/ebreak.S",
  "rv64i_m/privilege/src/ecall.S",
  "rv64i_m/privilege/src/misalign2-jalr-01.S",
  "rv64i_m/privilege/src/misalign-beq-01.S",
  "rv64i_m/privilege/src/misalign-bge-01.S",
  "rv64i_m/privilege/src/misalign-bgeu-01.S",
  "rv64i_m/privilege/src/misalign-blt-01.S",
  "rv64i_m/privilege/src/misalign-bltu-01.S",
  "rv64i_m/privilege/src/misalign-bne-01.S",
  "rv64i_m/privilege/src/misalign-jal-01.S",
  "rv64i_m/privilege/src/misalign-ld-01.S",
  "rv64i_m/privilege/src/misalign-lh-01.S",
  "rv64i_m/privilege/src/misalign-lhu-01.S",
  "rv64i_m/privilege/src/misalign-lw-01.S",
  "rv64i_m/privilege/src/misalign-lwu-01.S",
  "rv64i_m/privilege/src/misalign-sd-01.S",
  "rv64i_m/privilege/src/misalign-sh-01.S",
  "rv64i_m/privilege/src/misalign-sw-01.S"
};

string arch64zifencei[] = '{
  `RISCVARCHTEST,
  "rv64i_m/Zifencei/src/Fencei.S"
};

string arch64zicond[] = '{
  `RISCVARCHTEST,
  "rv64i_m/Zicond/src/czero.eqz-01.S",
  "rv64i_m/Zicond/src/czero.nez-01.S"
};

string arch32a_amo[] = '{
  `RISCVARCHTEST,
  "rv32i_m/A/src/amoadd.w-01.S",
  "rv32i_m/A/src/amoand.w-01.S",
  "rv32i_m/A/src/amomax.w-01.S",
  "rv32i_m/A/src/amomaxu.w-01.S",
  "rv32i_m/A/src/amomin.w-01.S",
  "rv32i_m/A/src/amominu.w-01.S",
  "rv32i_m/A/src/amoor.w-01.S",
  "rv32i_m/A/src/amoswap.w-01.S",
  "rv32i_m/A/src/amoxor.w-01.S"
};


string arch32zifencei[] = '{
  `RISCVARCHTEST,
  "rv32i_m/Zifencei/src/Fencei.S"
};

string arch32zicond[] = '{
  `RISCVARCHTEST,
  "rv32i_m/Zicond/src/czero.eqz-01.S",
  "rv32i_m/Zicond/src/czero.nez-01.S"
};

string arch32zba[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/sh1add-01.S",
  "rv32i_m/B/src/sh2add-01.S",
  "rv32i_m/B/src/sh3add-01.S"
};

string arch32zbb[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/max-01.S",
  "rv32i_m/B/src/maxu-01.S",
  "rv32i_m/B/src/min-01.S",
  "rv32i_m/B/src/minu-01.S",
  "rv32i_m/B/src/orcb_32-01.S",
  "rv32i_m/B/src/rev8_32-01.S",
  "rv32i_m/B/src/andn-01.S",
  "rv32i_m/B/src/orn-01.S",
  "rv32i_m/B/src/xnor-01.S",
  "rv32i_m/B/src/zext.h_32-01.S",
  "rv32i_m/B/src/sext.b-01.S",
  "rv32i_m/B/src/sext.h-01.S",
  "rv32i_m/B/src/clz-01.S",
  "rv32i_m/B/src/cpop-01.S",
  "rv32i_m/B/src/ctz-01.S",
  "rv32i_m/B/src/ror-01.S",
  "rv32i_m/B/src/rori-01.S",
  "rv32i_m/B/src/rol-01.S"
};

string arch32zbc[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/clmul-01.S",
  "rv32i_m/B/src/clmulh-01.S",
  "rv32i_m/B/src/clmulr-01.S"
};

string arch32zbs[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/bclr-01.S",
  "rv32i_m/B/src/bclri-01.S",
  "rv32i_m/B/src/bext-01.S",
  "rv32i_m/B/src/bexti-01.S",
  "rv32i_m/B/src/binv-01.S",
  "rv32i_m/B/src/binvi-01.S",
  "rv32i_m/B/src/bset-01.S",
  "rv32i_m/B/src/bseti-01.S"
};

string arch32zbkc[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/clmul-01.S",
  "rv32i_m/B/src/clmulh-01.S"
};

string arch32zbkx[] = '{
  `RISCVARCHTEST,
  "rv32i_m/K/src/xperm8-01.S",
  "rv32i_m/K/src/xperm4-01.S"
};

string arch32zknd[] = '{
  `RISCVARCHTEST,
  "rv32i_m/K/src/aes32dsi-01.S",
  "rv32i_m/K/src/aes32dsmi-01.S"
};

string arch32zkne[] = '{
  `RISCVARCHTEST,
  "rv32i_m/K/src/aes32esi-01.S",
  "rv32i_m/K/src/aes32esmi-01.S"
};

string arch32zknh[] = '{
  `RISCVARCHTEST,
  "rv32i_m/K/src/sha256sig0-01.S",
  "rv32i_m/K/src/sha256sig1-01.S",
  "rv32i_m/K/src/sha256sum0-01.S",
  "rv32i_m/K/src/sha256sum1-01.S",
  "rv32i_m/K/src/sha512sig0h-01.S",
  "rv32i_m/K/src/sha512sig0l-01.S",
  "rv32i_m/K/src/sha512sig1h-01.S",
  "rv32i_m/K/src/sha512sig1l-01.S",
  "rv32i_m/K/src/sha512sum0r-01.S",
  "rv32i_m/K/src/sha512sum1r-01.S"
};

string arch32zbkb[] = '{
  `RISCVARCHTEST,
  "rv32i_m/B/src/ror-01.S",
  "rv32i_m/B/src/rol-01.S",
  "rv32i_m/B/src/rori-01.S",
  "rv32i_m/B/src/andn-01.S",
  "rv32i_m/B/src/orn-01.S",
  "rv32i_m/B/src/xnor-01.S",
  "rv32i_m/B/src/rev8_32-01.S",
  "rv32i_m/K/src/pack-01.S",
  "rv32i_m/K/src/packh-01.S",
  "rv32i_m/K/src/brev8_32-01.S",
  "rv32i_m/K/src/zip-01.S",
  "rv32i_m/K/src/unzip-01.S"
};

string arch64zbkb[] = '{
  `RISCVARCHTEST,
  "rv64i_m/B/src/ror-01.S",
  "rv64i_m/B/src/rol-01.S",
  "rv64i_m/B/src/rori-01.S",
  "rv64i_m/B/src/rorw-01.S",
  "rv64i_m/B/src/rolw-01.S",
  "rv64i_m/B/src/roriw-01.S",
  "rv64i_m/B/src/andn-01.S",
  "rv64i_m/B/src/orn-01.S",
  "rv64i_m/B/src/xnor-01.S",
  "rv64i_m/B/src/rev8-01.S",
  "rv64i_m/K/src/pack-01.S",
  "rv64i_m/K/src/packh-01.S",
  "rv64i_m/K/src/packw-01.S",
  "rv64i_m/K/src/brev8-01.S"
};

string arch64m[] = '{
  `RISCVARCHTEST,
  "rv64i_m/M/src/div-01.S",
  "rv64i_m/M/src/divu-01.S",
  "rv64i_m/M/src/divuw-01.S",
  "rv64i_m/M/src/divw-01.S",
  "rv64i_m/M/src/mul-01.S",
  "rv64i_m/M/src/mulh-01.S",
  "rv64i_m/M/src/mulhsu-01.S",
  "rv64i_m/M/src/mulhu-01.S",
  "rv64i_m/M/src/mulw-01.S",
  "rv64i_m/M/src/rem-01.S",
  "rv64i_m/M/src/remu-01.S",
  "rv64i_m/M/src/remuw-01.S",
  "rv64i_m/M/src/remw-01.S"
};

string arch64a_amo[] = '{
  `RISCVARCHTEST,
  "rv64i_m/A/src/amoadd.w-01.S",
  "rv64i_m/A/src/amoand.w-01.S",
  "rv64i_m/A/src/amomax.w-01.S",
  "rv64i_m/A/src/amomaxu.w-01.S",
  "rv64i_m/A/src/amomin.w-01.S",
  "rv64i_m/A/src/amominu.w-01.S",
  "rv64i_m/A/src/amoor.w-01.S",
  "rv64i_m/A/src/amoswap.w-01.S",
  "rv64i_m/A/src/amoxor.w-01.S",
  "rv64i_m/A/src/amoadd.d-01.S",
  "rv64i_m/A/src/amoand.d-01.S",
  "rv64i_m/A/src/amomax.d-01.S",
  "rv64i_m/A/src/amomaxu.d-01.S",
  "rv64i_m/A/src/amomin.d-01.S",
  "rv64i_m/A/src/amominu.d-01.S",
  "rv64i_m/A/src/amoor.d-01.S",
  "rv64i_m/A/src/amoswap.d-01.S",
  "rv64i_m/A/src/amoxor.d-01.S"
};

string arch64c[] = '{
  `RISCVARCHTEST,
  "rv64i_m/C/src/cadd-01.S",
  "rv64i_m/C/src/caddi-01.S",
  "rv64i_m/C/src/caddi16sp-01.S",
  "rv64i_m/C/src/caddi4spn-01.S",
  "rv64i_m/C/src/caddiw-01.S",
  "rv64i_m/C/src/caddw-01.S",
  "rv64i_m/C/src/cand-01.S",
  "rv64i_m/C/src/candi-01.S",
  "rv64i_m/C/src/cbeqz-01.S",
  "rv64i_m/C/src/cbnez-01.S",
  "rv64i_m/C/src/cj-01.S",
  "rv64i_m/C/src/cjalr-01.S",
  "rv64i_m/C/src/cjr-01.S",
  "rv64i_m/C/src/cld-01.S",
  "rv64i_m/C/src/cldsp-01.S",
  "rv64i_m/C/src/cli-01.S",
  "rv64i_m/C/src/clui-01.S",
  "rv64i_m/C/src/clw-01.S",
  "rv64i_m/C/src/clwsp-01.S",
  "rv64i_m/C/src/cmv-01.S",
  "rv64i_m/C/src/cnop-01.S",
  "rv64i_m/C/src/cor-01.S",
  "rv64i_m/C/src/csd-01.S",
  "rv64i_m/C/src/csdsp-01.S",
  "rv64i_m/C/src/cslli-01.S",
  "rv64i_m/C/src/csrai-01.S",
  "rv64i_m/C/src/csrli-01.S",
  "rv64i_m/C/src/csub-01.S",
  "rv64i_m/C/src/csubw-01.S",
  "rv64i_m/C/src/csw-01.S",
  "rv64i_m/C/src/cswsp-01.S",
  "rv64i_m/C/src/cxor-01.S"
  //"rv64i_m/C/src/misalign1-cjalr-01.S", // no longer in repo
  //"rv64i_m/C/src/misalign1-cjr-01.S"
};

string arch64cpriv[] = '{
  // `RISCVARCHTEST,
  "rv64i_m/C/src/cebreak-01.S"
};

string arch64zcd[] = '{
  // `RISCVARCHTEST,
  "rv64i_m/D_Zcd/src/c.fld-01.S",
  "rv64i_m/D_Zcd/src/c.fldsp-01.S",
  "rv64i_m/D_Zcd/src/c.fsd-01.S",
  "rv64i_m/D_Zcd/src/c.fsdsp-01.S"
};

string arch64i[] = '{
  `RISCVARCHTEST,
  "rv64i_m/I/src/add-01.S",
  "rv64i_m/I/src/addi-01.S",
  "rv64i_m/I/src/addiw-01.S",
  "rv64i_m/I/src/addw-01.S",
  "rv64i_m/I/src/and-01.S",
  "rv64i_m/I/src/andi-01.S",
  "rv64i_m/I/src/auipc-01.S",
  "rv64i_m/I/src/beq-01.S",
  "rv64i_m/I/src/bge-01.S",
  "rv64i_m/I/src/bgeu-01.S",
  "rv64i_m/I/src/blt-01.S",
  "rv64i_m/I/src/bltu-01.S",
  "rv64i_m/I/src/bne-01.S",
  "rv64i_m/I/src/fence-01.S",
  "rv64i_m/I/src/jal-01.S",
  "rv64i_m/I/src/jalr-01.S",
  "rv64i_m/I/src/lb-align-01.S",
  "rv64i_m/I/src/lbu-align-01.S",
  "rv64i_m/I/src/ld-align-01.S",
  "rv64i_m/I/src/lh-align-01.S",
  "rv64i_m/I/src/lhu-align-01.S",
  "rv64i_m/I/src/lui-01.S",
  "rv64i_m/I/src/lw-align-01.S",
  "rv64i_m/I/src/lwu-align-01.S",
  "rv64i_m/I/src/or-01.S",
  "rv64i_m/I/src/ori-01.S",
  "rv64i_m/I/src/sb-align-01.S",
  "rv64i_m/I/src/sd-align-01.S",
  "rv64i_m/I/src/sh-align-01.S",
  "rv64i_m/I/src/sll-01.S",
  "rv64i_m/I/src/slli-01.S",
  "rv64i_m/I/src/slliw-01.S",
  "rv64i_m/I/src/sllw-01.S",
  "rv64i_m/I/src/slt-01.S",
  "rv64i_m/I/src/slti-01.S",
  "rv64i_m/I/src/sltiu-01.S",
  "rv64i_m/I/src/sltu-01.S",
  "rv64i_m/I/src/sra-01.S",
  "rv64i_m/I/src/srai-01.S",
  "rv64i_m/I/src/sraiw-01.S",
  "rv64i_m/I/src/sraw-01.S",
  "rv64i_m/I/src/srl-01.S",
  "rv64i_m/I/src/srli-01.S",
  "rv64i_m/I/src/srliw-01.S",
  "rv64i_m/I/src/srlw-01.S",
  "rv64i_m/I/src/sub-01.S",
  "rv64i_m/I/src/subw-01.S",
  "rv64i_m/I/src/sw-align-01.S",
  "rv64i_m/I/src/xor-01.S",
  "rv64i_m/I/src/xori-01.S"
};

string arch64f_fma[] = '{
  `RISCVARCHTEST,
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-001.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-002.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-003.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-004.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-005.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-006.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-007.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-008.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-009.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-010.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-011.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-012.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-013.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-014.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-015.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-016.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-017.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-018.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-019.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-020.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-021.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-022.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-023.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-024.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-025.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-026.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-027.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-028.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-029.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-030.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-031.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-032.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-033.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-034.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-035.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-036.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-037.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-038.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-039.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-040.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-041.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-042.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-043.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-044.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-045.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-046.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-047.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-048.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-049.S",
  // "rv64i_m/F/src/fmadd_b15/fmadd_b15-050.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-001.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-002.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-003.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-004.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-005.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-006.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-007.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-008.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-009.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-010.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-011.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-012.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-013.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-014.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-015.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-016.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-017.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-018.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-019.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-020.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-021.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-022.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-023.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-024.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-025.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-026.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-027.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-028.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-029.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-030.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-031.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-032.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-033.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-034.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-035.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-036.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-037.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-038.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-039.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-040.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-041.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-042.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-043.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-044.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-045.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-046.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-047.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-048.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-049.S",
  "rv64i_m/F/src/fmsub_b15/fmsub_b15-050.S"
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-001.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-002.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-003.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-004.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-005.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-006.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-007.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-008.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-009.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-010.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-011.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-012.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-013.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-014.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-015.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-016.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-017.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-018.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-019.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-020.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-021.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-022.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-023.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-024.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-025.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-026.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-027.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-028.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-029.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-030.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-031.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-032.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-033.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-034.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-035.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-036.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-037.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-038.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-039.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-040.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-041.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-042.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-043.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-044.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-045.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-046.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-047.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-048.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-049.S",
  // "rv64i_m/F/src/fnmadd_b15/fnmadd_b15-050.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-001.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-002.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-003.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-004.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-005.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-006.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-007.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-008.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-009.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-010.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-011.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-012.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-013.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-014.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-015.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-016.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-017.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-018.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-019.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-020.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-021.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-022.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-023.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-024.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-025.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-026.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-027.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-028.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-029.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-030.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-031.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-032.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-033.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-034.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-035.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-036.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-037.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-038.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-039.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-040.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-041.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-042.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-043.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-044.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-045.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-046.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-047.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-048.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-049.S",
  // "rv64i_m/F/src/fnmsub_b15/fnmsub_b15-050.S"
};

string arch64zfh_fma[] = '{
  `RISCVARCHTEST,
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-001.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-002.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-003.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-004.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-005.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-006.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-007.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-008.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-009.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-010.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-011.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-012.S",
  "rv64i_m/Zfh/src/fmadd_b15/fmadd_b15-013.S",

  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-001.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-002.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-003.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-004.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-005.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-006.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-007.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-008.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-009.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-010.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-011.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-012.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-013.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-014.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-015.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-016.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-017.S",
  "rv64i_m/Zfh/src/fmadd_b1/fmadd_b1-018.S",

  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-001.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-002.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-003.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-004.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-005.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-006.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-007.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-008.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-009.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-010.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-011.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-012.S",
  "rv64i_m/Zfh/src/fmsub_b15/fmsub_b15-013.S",

  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-001.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-002.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-003.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-004.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-005.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-006.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-007.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-008.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-009.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-010.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-011.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-012.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-013.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-014.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-015.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-016.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-017.S",
  "rv64i_m/Zfh/src/fmsub_b1/fmsub_b1-018.S",

  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-001.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-002.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-003.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-004.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-005.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-006.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-007.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-008.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-009.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-010.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-011.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-012.S",
  "rv64i_m/Zfh/src/fnmadd_b15/fnmadd_b15-013.S",

  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-001.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-002.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-003.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-004.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-005.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-006.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-007.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-008.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-009.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-010.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-011.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-012.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-013.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-014.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-015.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-016.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-017.S",
  "rv64i_m/Zfh/src/fnmadd_b1/fnmadd_b1-018.S",

  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-001.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-002.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-003.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-004.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-005.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-006.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-007.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-008.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-009.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-010.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-011.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-012.S",
  "rv64i_m/Zfh/src/fnmsub_b15/fnmsub_b15-013.S",

  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-001.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-002.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-003.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-004.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-005.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-006.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-007.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-008.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-009.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-010.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-011.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-012.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-013.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-014.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-015.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-016.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-017.S",
  "rv64i_m/Zfh/src/fnmsub_b1/fnmsub_b1-018.S"
};

string arch64f_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv64i_m/F/src/fdiv_b20-01.S",
  "rv64i_m/F/src/fdiv_b1-01.S",
  "rv64i_m/F/src/fdiv_b2-01.S",
  "rv64i_m/F/src/fdiv_b21-01.S",
  "rv64i_m/F/src/fdiv_b3-01.S",
  "rv64i_m/F/src/fdiv_b4-01.S",
  "rv64i_m/F/src/fdiv_b5-01.S",
  "rv64i_m/F/src/fdiv_b6-01.S",
  "rv64i_m/F/src/fdiv_b7-01.S",
  "rv64i_m/F/src/fdiv_b8-01.S",
  "rv64i_m/F/src/fdiv_b9-01.S",
  "rv64i_m/F/src/fsqrt_b1-01.S",
  "rv64i_m/F/src/fsqrt_b20-01.S",
  "rv64i_m/F/src/fsqrt_b2-01.S",
  "rv64i_m/F/src/fsqrt_b3-01.S",
  "rv64i_m/F/src/fsqrt_b4-01.S",
  "rv64i_m/F/src/fsqrt_b5-01.S",
  "rv64i_m/F/src/fsqrt_b7-01.S",
  "rv64i_m/F/src/fsqrt_b8-01.S",
  "rv64i_m/F/src/fsqrt_b9-01.S"
};

string arch64f[] = '{
  `RISCVARCHTEST,
  "rv64i_m/F/src/fadd_b10-01.S",
  "rv64i_m/F/src/fadd_b1-01.S",
  "rv64i_m/F/src/fadd_b11-01.S",
  "rv64i_m/F/src/fadd_b12-01.S",
  "rv64i_m/F/src/fadd_b13-01.S",
  "rv64i_m/F/src/fadd_b2-01.S",
  "rv64i_m/F/src/fadd_b3-01.S",
  "rv64i_m/F/src/fadd_b4-01.S",
  "rv64i_m/F/src/fadd_b5-01.S",
  "rv64i_m/F/src/fadd_b7-01.S",
  "rv64i_m/F/src/fadd_b8-01.S",
  "rv64i_m/F/src/fclass_b1-01.S",
  "rv64i_m/F/src/fcvt.s.l_b25-01.S",
  "rv64i_m/F/src/fcvt.s.l_b26-01.S",
  "rv64i_m/F/src/fcvt.s.lu_b25-01.S",
  "rv64i_m/F/src/fcvt.s.lu_b26-01.S",
  "rv64i_m/F/src/fcvt.l.s_b1-01.S",
  "rv64i_m/F/src/fcvt.l.s_b22-01.S",
  "rv64i_m/F/src/fcvt.l.s_b23-01.S",
  "rv64i_m/F/src/fcvt.l.s_b24-01.S",
  "rv64i_m/F/src/fcvt.l.s_b27-01.S",
  "rv64i_m/F/src/fcvt.l.s_b28-01.S",
  "rv64i_m/F/src/fcvt.l.s_b29-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b1-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b22-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b23-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b24-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b27-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b28-01.S",
  "rv64i_m/F/src/fcvt.lu.s_b29-01.S",
  "rv64i_m/F/src/fcvt.s.w_b25-01.S",
  "rv64i_m/F/src/fcvt.s.w_b26-01.S",
  "rv64i_m/F/src/fcvt.s.wu_b25-01.S",
  "rv64i_m/F/src/fcvt.s.wu_b26-01.S",
  "rv64i_m/F/src/fcvt.w.s_b1-01.S",
  "rv64i_m/F/src/fcvt.w.s_b22-01.S",
  "rv64i_m/F/src/fcvt.w.s_b23-01.S",
  "rv64i_m/F/src/fcvt.w.s_b24-01.S",
  "rv64i_m/F/src/fcvt.w.s_b27-01.S",
  "rv64i_m/F/src/fcvt.w.s_b28-01.S",
  "rv64i_m/F/src/fcvt.w.s_b29-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b1-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b22-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b23-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b24-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b27-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b28-01.S",
  "rv64i_m/F/src/fcvt.wu.s_b29-01.S",
  "rv64i_m/F/src/feq_b1-01.S",
  "rv64i_m/F/src/feq_b19-01.S",
  "rv64i_m/F/src/fle_b1-01.S",
  "rv64i_m/F/src/fle_b19-01.S",
  "rv64i_m/F/src/flt_b1-01.S",
  "rv64i_m/F/src/flt_b19-01.S",
  "rv64i_m/F/src/flw-align-01.S",
  //"rv64i_m/F/src/fmadd_b1-01.S",
  "rv64i_m/F/src/fmadd_b14-01.S",
  "rv64i_m/F/src/fmadd_b16-01.S",
  "rv64i_m/F/src/fmadd_b17-01.S",
  "rv64i_m/F/src/fmadd_b18-01.S",
  "rv64i_m/F/src/fmadd_b2-01.S",
  "rv64i_m/F/src/fmadd_b3-01.S",
  "rv64i_m/F/src/fmadd_b4-01.S",
  "rv64i_m/F/src/fmadd_b5-01.S",
  "rv64i_m/F/src/fmadd_b6-01.S",
  "rv64i_m/F/src/fmadd_b7-01.S",
  "rv64i_m/F/src/fmadd_b8-01.S",
  "rv64i_m/F/src/fmax_b1-01.S",
  "rv64i_m/F/src/fmax_b19-01.S",
  "rv64i_m/F/src/fmin_b1-01.S",
  "rv64i_m/F/src/fmin_b19-01.S",
  "rv64i_m/F/src/fmsub_b1-01.S",
  "rv64i_m/F/src/fmsub_b14-01.S",
  "rv64i_m/F/src/fmsub_b16-01.S",
  "rv64i_m/F/src/fmsub_b17-01.S",
  "rv64i_m/F/src/fmsub_b18-01.S",
  "rv64i_m/F/src/fmsub_b2-01.S",
  "rv64i_m/F/src/fmsub_b3-01.S",
  "rv64i_m/F/src/fmsub_b4-01.S",
  "rv64i_m/F/src/fmsub_b5-01.S",
  "rv64i_m/F/src/fmsub_b6-01.S",
  "rv64i_m/F/src/fmsub_b7-01.S",
  "rv64i_m/F/src/fmsub_b8-01.S",
  "rv64i_m/F/src/fmul_b1-01.S",
  "rv64i_m/F/src/fmul_b2-01.S",
  "rv64i_m/F/src/fmul_b3-01.S",
  "rv64i_m/F/src/fmul_b4-01.S",
  "rv64i_m/F/src/fmul_b5-01.S",
  "rv64i_m/F/src/fmul_b6-01.S",
  "rv64i_m/F/src/fmul_b7-01.S",
  "rv64i_m/F/src/fmul_b8-01.S",
  "rv64i_m/F/src/fmul_b9-01.S",
  "rv64i_m/F/src/fmv.w.x_b25-01.S",
  "rv64i_m/F/src/fmv.w.x_b26-01.S",
  "rv64i_m/F/src/fmv.x.w_b1-01.S",
  "rv64i_m/F/src/fmv.x.w_b22-01.S",
  "rv64i_m/F/src/fmv.x.w_b23-01.S",
  "rv64i_m/F/src/fmv.x.w_b24-01.S",
  "rv64i_m/F/src/fmv.x.w_b27-01.S",
  "rv64i_m/F/src/fmv.x.w_b28-01.S",
  "rv64i_m/F/src/fmv.x.w_b29-01.S",
  "rv64i_m/F/src/fnmadd_b1-01.S",
  "rv64i_m/F/src/fnmadd_b14-01.S",
  "rv64i_m/F/src/fnmadd_b16-01.S",
  "rv64i_m/F/src/fnmadd_b17-01.S",
  "rv64i_m/F/src/fnmadd_b18-01.S",
  "rv64i_m/F/src/fnmadd_b2-01.S",
  "rv64i_m/F/src/fnmadd_b3-01.S",
  "rv64i_m/F/src/fnmadd_b4-01.S",
  "rv64i_m/F/src/fnmadd_b5-01.S",
  "rv64i_m/F/src/fnmadd_b6-01.S",
  "rv64i_m/F/src/fnmadd_b7-01.S",
  "rv64i_m/F/src/fnmadd_b8-01.S",
  "rv64i_m/F/src/fnmsub_b1-01.S",
  "rv64i_m/F/src/fnmsub_b14-01.S",
  "rv64i_m/F/src/fnmsub_b16-01.S",
  "rv64i_m/F/src/fnmsub_b17-01.S",
  "rv64i_m/F/src/fnmsub_b18-01.S",
  "rv64i_m/F/src/fnmsub_b2-01.S",
  "rv64i_m/F/src/fnmsub_b3-01.S",
  "rv64i_m/F/src/fnmsub_b4-01.S",
  "rv64i_m/F/src/fnmsub_b5-01.S",
  "rv64i_m/F/src/fnmsub_b6-01.S",
  "rv64i_m/F/src/fnmsub_b7-01.S",
  "rv64i_m/F/src/fnmsub_b8-01.S",
  "rv64i_m/F/src/fsgnj_b1-01.S",
  "rv64i_m/F/src/fsgnjn_b1-01.S",
  "rv64i_m/F/src/fsgnjx_b1-01.S",
  "rv64i_m/F/src/fsub_b10-01.S",
  "rv64i_m/F/src/fsub_b1-01.S",
  "rv64i_m/F/src/fsub_b11-01.S",
  "rv64i_m/F/src/fsub_b12-01.S",
  "rv64i_m/F/src/fsub_b13-01.S",
  "rv64i_m/F/src/fsub_b2-01.S",
  "rv64i_m/F/src/fsub_b3-01.S",
  "rv64i_m/F/src/fsub_b4-01.S",
  "rv64i_m/F/src/fsub_b5-01.S",
  "rv64i_m/F/src/fsub_b7-01.S",
  "rv64i_m/F/src/fsub_b8-01.S",
  "rv64i_m/F/src/fsw-align-01.S"
};

string arch64zfh_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv64i_m/Zfh/src/fdiv_b20-01.S",
  "rv64i_m/Zfh/src/fdiv_b1-01.S",
  "rv64i_m/Zfh/src/fdiv_b2-01.S",
  "rv64i_m/Zfh/src/fdiv_b21-01.S",
  "rv64i_m/Zfh/src/fdiv_b3-01.S",
  "rv64i_m/Zfh/src/fdiv_b4-01.S",
  "rv64i_m/Zfh/src/fdiv_b5-01.S",
  "rv64i_m/Zfh/src/fdiv_b6-01.S",
  "rv64i_m/Zfh/src/fdiv_b7-01.S",
  "rv64i_m/Zfh/src/fdiv_b8-01.S",
  "rv64i_m/Zfh/src/fdiv_b9-01.S",
  "rv64i_m/Zfh/src/fsqrt_b1-01.S",
  "rv64i_m/Zfh/src/fsqrt_b20-01.S",
  "rv64i_m/Zfh/src/fsqrt_b2-01.S",
  "rv64i_m/Zfh/src/fsqrt_b3-01.S",
  "rv64i_m/Zfh/src/fsqrt_b4-01.S",
  "rv64i_m/Zfh/src/fsqrt_b5-01.S",
  "rv64i_m/Zfh/src/fsqrt_b7-01.S",
  "rv64i_m/Zfh/src/fsqrt_b8-01.S",
  "rv64i_m/Zfh/src/fsqrt_b9-01.S"
};

string arch64zfh[] = '{
  `RISCVARCHTEST,
  "rv64i_m/Zfh/src/fadd_b10-01.S",
  "rv64i_m/Zfh/src/fadd_b1-01.S",
  "rv64i_m/Zfh/src/fadd_b11-01.S",
  "rv64i_m/Zfh/src/fadd_b12-01.S",
  "rv64i_m/Zfh/src/fadd_b13-01.S",
  "rv64i_m/Zfh/src/fadd_b2-01.S",
  "rv64i_m/Zfh/src/fadd_b3-01.S",
  "rv64i_m/Zfh/src/fadd_b4-01.S",
  "rv64i_m/Zfh/src/fadd_b5-01.S",
  "rv64i_m/Zfh/src/fadd_b7-01.S",
  "rv64i_m/Zfh/src/fadd_b8-01.S",
  "rv64i_m/Zfh/src/fclass_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.h.s_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.h.w_b25-01.S",
  "rv64i_m/Zfh/src/fcvt.h.w_b26-01.S",
  "rv64i_m/Zfh/src/fcvt.h.wu_b25-01.S",
  "rv64i_m/Zfh/src/fcvt.h.wu_b26-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.s.h_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.w.h_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.wu.h_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.h.l_b25-01.S",
  "rv64i_m/Zfh/src/fcvt.h.l_b26-01.S",
  "rv64i_m/Zfh/src/fcvt.h.lu_b25-01.S",
  "rv64i_m/Zfh/src/fcvt.h.lu_b26-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.l.h_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.lu.h_b29-01.S",
  "rv64i_m/Zfh/src/feq_b1-01.S",
  "rv64i_m/Zfh/src/feq_b19-01.S",
  "rv64i_m/Zfh/src/fle_b1-01.S",
  "rv64i_m/Zfh/src/fle_b19-01.S",
  "rv64i_m/Zfh/src/flt_b1-01.S",
  "rv64i_m/Zfh/src/flt_b19-01.S",
  "rv64i_m/Zfh/src/flh-align-01.S",
  "rv64i_m/Zfh/src/fmax_b1-01.S",
  "rv64i_m/Zfh/src/fmax_b19-01.S",
  "rv64i_m/Zfh/src/fmin_b1-01.S",
  "rv64i_m/Zfh/src/fmin_b19-01.S",
  "rv64i_m/Zfh/src/fmul_b1-01.S",
  "rv64i_m/Zfh/src/fmul_b2-01.S",
  "rv64i_m/Zfh/src/fmul_b3-01.S",
  "rv64i_m/Zfh/src/fmul_b4-01.S",
  "rv64i_m/Zfh/src/fmul_b5-01.S",
  "rv64i_m/Zfh/src/fmul_b6-01.S",
  "rv64i_m/Zfh/src/fmul_b7-01.S",
  "rv64i_m/Zfh/src/fmul_b8-01.S",
  "rv64i_m/Zfh/src/fmul_b9-01.S",
  "rv64i_m/Zfh/src/fmv.h.x_b25-01.S",
  "rv64i_m/Zfh/src/fmv.h.x_b26-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b1-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b22-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b23-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b24-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b27-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b28-01.S",
  "rv64i_m/Zfh/src/fmv.x.h_b29-01.S",
  "rv64i_m/Zfh/src/fsgnj_b1-01.S",
  "rv64i_m/Zfh/src/fsgnjn_b1-01.S",
  "rv64i_m/Zfh/src/fsgnjx_b1-01.S",
  "rv64i_m/Zfh/src/fsub_b10-01.S",
  "rv64i_m/Zfh/src/fsub_b1-01.S",
  "rv64i_m/Zfh/src/fsub_b11-01.S",
  "rv64i_m/Zfh/src/fsub_b12-01.S",
  "rv64i_m/Zfh/src/fsub_b13-01.S",
  "rv64i_m/Zfh/src/fsub_b2-01.S",
  "rv64i_m/Zfh/src/fsub_b3-01.S",
  "rv64i_m/Zfh/src/fsub_b4-01.S",
  "rv64i_m/Zfh/src/fsub_b5-01.S",
  "rv64i_m/Zfh/src/fsub_b7-01.S",
  "rv64i_m/Zfh/src/fsub_b8-01.S",
  "rv64i_m/Zfh/src/fsh-align-01.S",
  "rv64i_m/Zfh/src/fmadd_b14-01.S",
  "rv64i_m/Zfh/src/fmadd_b16-01.S",
  "rv64i_m/Zfh/src/fmadd_b17-01.S",
  "rv64i_m/Zfh/src/fmadd_b18-01.S",
  "rv64i_m/Zfh/src/fmadd_b2-01.S",
  "rv64i_m/Zfh/src/fmadd_b3-01.S",
  "rv64i_m/Zfh/src/fmadd_b4-01.S",
  "rv64i_m/Zfh/src/fmadd_b5-01.S",
  "rv64i_m/Zfh/src/fmadd_b6-01.S",
  "rv64i_m/Zfh/src/fmadd_b7-01.S",
  "rv64i_m/Zfh/src/fmadd_b8-01.S",
  "rv64i_m/Zfh/src/fmsub_b14-01.S",
  "rv64i_m/Zfh/src/fmsub_b16-01.S",
  "rv64i_m/Zfh/src/fmsub_b17-01.S",
  "rv64i_m/Zfh/src/fmsub_b18-01.S",
  "rv64i_m/Zfh/src/fmsub_b2-01.S",
  "rv64i_m/Zfh/src/fmsub_b3-01.S",
  "rv64i_m/Zfh/src/fmsub_b4-01.S",
  "rv64i_m/Zfh/src/fmsub_b5-01.S",
  "rv64i_m/Zfh/src/fmsub_b6-01.S",
  "rv64i_m/Zfh/src/fmsub_b7-01.S",
  "rv64i_m/Zfh/src/fmsub_b8-01.S",
  "rv64i_m/Zfh/src/fnmadd_b14-01.S",
  "rv64i_m/Zfh/src/fnmadd_b16-01.S",
  "rv64i_m/Zfh/src/fnmadd_b17-01.S",
  "rv64i_m/Zfh/src/fnmadd_b18-01.S",
  "rv64i_m/Zfh/src/fnmadd_b2-01.S",
  "rv64i_m/Zfh/src/fnmadd_b3-01.S",
  "rv64i_m/Zfh/src/fnmadd_b4-01.S",
  "rv64i_m/Zfh/src/fnmadd_b5-01.S",
  "rv64i_m/Zfh/src/fnmadd_b6-01.S",
  "rv64i_m/Zfh/src/fnmadd_b7-01.S",
  "rv64i_m/Zfh/src/fnmadd_b8-01.S",
  "rv64i_m/Zfh/src/fnmsub_b14-01.S",
  "rv64i_m/Zfh/src/fnmsub_b16-01.S",
  "rv64i_m/Zfh/src/fnmsub_b17-01.S",
  "rv64i_m/Zfh/src/fnmsub_b18-01.S",
  "rv64i_m/Zfh/src/fnmsub_b2-01.S",
  "rv64i_m/Zfh/src/fnmsub_b3-01.S",
  "rv64i_m/Zfh/src/fnmsub_b4-01.S",
  "rv64i_m/Zfh/src/fnmsub_b5-01.S",
  "rv64i_m/Zfh/src/fnmsub_b6-01.S",
  "rv64i_m/Zfh/src/fnmsub_b7-01.S",
  "rv64i_m/Zfh/src/fnmsub_b8-01.S"
};

string arch64zfh_d[] = '{
  // `RISCVARCHTEST,
  "rv64i_m/Zfh/src/fcvt.d.h_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.d.h_b29-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b1-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b22-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b23-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b24-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b27-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b28-01.S",
  "rv64i_m/Zfh/src/fcvt.h.d_b29-01.S"
};

string arch64d_fma[] = '{
  `RISCVARCHTEST,
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-001.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-002.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-003.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-004.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-005.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-006.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-007.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-008.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-009.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-010.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-011.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-012.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-013.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-014.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-015.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-016.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-017.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-018.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-019.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-020.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-021.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-022.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-023.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-024.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-025.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-026.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-027.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-028.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-029.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-030.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-031.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-032.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-033.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-034.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-035.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-036.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-037.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-038.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-039.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-040.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-041.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-042.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-043.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-044.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-045.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-046.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-047.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-048.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-049.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-050.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-051.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-052.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-053.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-054.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-055.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-056.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-057.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-058.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-059.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-060.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-061.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-062.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-063.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-064.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-065.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-066.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-067.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-068.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-069.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-070.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-071.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-072.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-073.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-074.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-075.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-076.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-077.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-078.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-079.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-080.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-081.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-082.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-083.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-084.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-085.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-086.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-087.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-088.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-089.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-090.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-091.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-092.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-093.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-094.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-095.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-096.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-097.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-098.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-099.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-100.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-101.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-102.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-103.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-104.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-105.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-106.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-107.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-108.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-109.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-110.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-111.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-112.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-113.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-114.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-115.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-116.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-117.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-118.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-119.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-120.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-121.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-122.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-123.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-124.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-125.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-126.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-127.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-128.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-129.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-130.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-131.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-132.S",
  // "rv64i_m/D/src/fmadd.d_b15/fmadd.d_b15-133.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-001.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-002.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-003.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-004.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-005.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-006.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-007.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-008.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-009.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-010.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-011.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-012.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-013.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-014.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-015.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-016.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-017.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-018.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-019.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-020.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-021.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-022.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-023.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-024.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-025.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-026.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-027.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-028.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-029.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-030.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-031.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-032.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-033.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-034.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-035.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-036.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-037.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-038.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-039.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-040.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-041.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-042.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-043.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-044.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-045.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-046.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-047.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-048.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-049.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-050.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-051.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-052.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-053.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-054.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-055.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-056.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-057.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-058.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-059.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-060.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-061.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-062.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-063.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-064.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-065.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-066.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-067.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-068.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-069.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-070.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-071.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-072.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-073.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-074.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-075.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-076.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-077.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-078.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-079.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-080.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-081.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-082.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-083.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-084.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-085.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-086.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-087.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-088.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-089.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-090.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-091.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-092.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-093.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-094.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-095.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-096.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-097.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-098.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-099.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-100.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-101.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-102.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-103.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-104.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-105.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-106.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-107.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-108.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-109.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-110.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-111.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-112.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-113.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-114.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-115.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-116.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-117.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-118.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-119.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-120.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-121.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-122.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-123.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-124.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-125.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-126.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-127.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-128.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-129.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-130.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-131.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-132.S",
  // "rv64i_m/D/src/fmsub.d_b15/fmsub.d_b15-133.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-001.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-002.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-003.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-004.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-005.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-006.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-007.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-008.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-009.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-010.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-011.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-012.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-013.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-014.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-015.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-016.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-017.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-018.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-019.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-020.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-021.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-022.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-023.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-024.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-025.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-026.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-027.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-028.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-029.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-030.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-031.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-032.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-033.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-034.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-035.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-036.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-037.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-038.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-039.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-040.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-041.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-042.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-043.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-044.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-045.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-046.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-047.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-048.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-049.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-050.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-051.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-052.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-053.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-054.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-055.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-056.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-057.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-058.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-059.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-060.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-061.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-062.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-063.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-064.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-065.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-066.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-067.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-068.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-069.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-070.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-071.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-072.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-073.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-074.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-075.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-076.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-077.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-078.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-079.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-080.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-081.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-082.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-083.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-084.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-085.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-086.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-087.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-088.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-089.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-090.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-091.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-092.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-093.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-094.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-095.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-096.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-097.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-098.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-099.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-100.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-101.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-102.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-103.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-104.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-105.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-106.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-107.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-108.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-109.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-110.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-111.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-112.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-113.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-114.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-115.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-116.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-117.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-118.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-119.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-120.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-121.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-122.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-123.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-124.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-125.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-126.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-127.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-128.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-129.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-130.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-131.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-132.S",
  "rv64i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-133.S"
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-001.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-002.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-003.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-004.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-005.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-006.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-007.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-008.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-009.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-010.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-011.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-012.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-013.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-014.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-015.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-016.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-017.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-018.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-019.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-020.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-021.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-022.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-023.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-024.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-025.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-026.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-027.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-028.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-029.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-030.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-031.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-032.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-033.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-034.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-035.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-036.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-037.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-038.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-039.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-040.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-041.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-042.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-043.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-044.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-045.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-046.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-047.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-048.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-049.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-050.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-051.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-052.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-053.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-054.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-055.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-056.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-057.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-058.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-059.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-060.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-061.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-062.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-063.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-064.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-065.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-066.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-067.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-068.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-069.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-070.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-071.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-072.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-073.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-074.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-075.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-076.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-077.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-078.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-079.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-080.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-081.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-082.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-083.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-084.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-085.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-086.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-087.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-088.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-089.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-090.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-091.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-092.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-093.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-094.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-095.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-096.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-097.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-098.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-099.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-100.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-101.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-102.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-103.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-104.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-105.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-106.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-107.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-108.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-109.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-110.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-111.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-112.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-113.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-114.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-115.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-116.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-117.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-118.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-119.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-120.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-121.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-122.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-123.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-124.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-125.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-126.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-127.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-128.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-129.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-130.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-131.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-132.S",
  // "rv64i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-133.S"
};

string arch64d_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv64i_m/D/src/fdiv.d_b1-01.S",
  "rv64i_m/D/src/fdiv.d_b20-01.S",
  "rv64i_m/D/src/fdiv.d_b2-01.S",
  "rv64i_m/D/src/fdiv.d_b21-01.S",
  "rv64i_m/D/src/fdiv.d_b3-01.S",
  "rv64i_m/D/src/fdiv.d_b4-01.S",
  "rv64i_m/D/src/fdiv.d_b5-01.S",
  "rv64i_m/D/src/fdiv.d_b6-01.S",
  "rv64i_m/D/src/fdiv.d_b7-01.S",
  "rv64i_m/D/src/fdiv.d_b8-01.S",
  "rv64i_m/D/src/fdiv.d_b9-01.S",
  "rv64i_m/D/src/fsqrt.d_b1-01.S",
  "rv64i_m/D/src/fsqrt.d_b20-01.S",
  "rv64i_m/D/src/fsqrt.d_b2-01.S",
  "rv64i_m/D/src/fsqrt.d_b3-01.S",
  "rv64i_m/D/src/fsqrt.d_b4-01.S",
  "rv64i_m/D/src/fsqrt.d_b5-01.S",
  "rv64i_m/D/src/fsqrt.d_b7-01.S",
  "rv64i_m/D/src/fsqrt.d_b8-01.S",
  "rv64i_m/D/src/fsqrt.d_b9-01.S"
};

string arch64d[] = '{
  `RISCVARCHTEST,
  // for speed
  "rv64i_m/D/src/fadd.d_b10-01.S",
  "rv64i_m/D/src/fadd.d_b1-01.S",
  "rv64i_m/D/src/fadd.d_b11-01.S",
  "rv64i_m/D/src/fadd.d_b12-01.S",
  "rv64i_m/D/src/fadd.d_b13-01.S",
  "rv64i_m/D/src/fadd.d_b2-01.S",
  "rv64i_m/D/src/fadd.d_b3-01.S",
  "rv64i_m/D/src/fadd.d_b4-01.S",
  "rv64i_m/D/src/fadd.d_b5-01.S",
  "rv64i_m/D/src/fadd.d_b7-01.S",
  "rv64i_m/D/src/fadd.d_b8-01.S",
  "rv64i_m/D/src/fclass.d_b1-01.S",
  "rv64i_m/D/src/fcvt.d.l_b25-01.S",
  "rv64i_m/D/src/fcvt.d.l_b26-01.S",
  "rv64i_m/D/src/fcvt.d.lu_b25-01.S",
  "rv64i_m/D/src/fcvt.d.lu_b26-01.S",
  "rv64i_m/D/src/fcvt.d.s_b1-01.S",
  "rv64i_m/D/src/fcvt.d.s_b22-01.S",
  "rv64i_m/D/src/fcvt.d.s_b23-01.S",
  "rv64i_m/D/src/fcvt.d.s_b24-01.S",
  "rv64i_m/D/src/fcvt.d.s_b27-01.S",
  "rv64i_m/D/src/fcvt.d.s_b28-01.S",
  "rv64i_m/D/src/fcvt.d.s_b29-01.S",
  "rv64i_m/D/src/fcvt.d.w_b25-01.S",
  "rv64i_m/D/src/fcvt.d.w_b26-01.S",
  "rv64i_m/D/src/fcvt.d.wu_b25-01.S",
  "rv64i_m/D/src/fcvt.d.wu_b26-01.S",
  "rv64i_m/D/src/fcvt.l.d_b1-01.S",
  "rv64i_m/D/src/fcvt.l.d_b22-01.S",
  "rv64i_m/D/src/fcvt.l.d_b23-01.S",
  "rv64i_m/D/src/fcvt.l.d_b24-01.S",
  "rv64i_m/D/src/fcvt.l.d_b27-01.S",
  "rv64i_m/D/src/fcvt.l.d_b28-01.S",
  "rv64i_m/D/src/fcvt.l.d_b29-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b1-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b22-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b23-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b24-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b27-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b28-01.S",
  "rv64i_m/D/src/fcvt.lu.d_b29-01.S",
  "rv64i_m/D/src/fcvt.s.d_b1-01.S",
  "rv64i_m/D/src/fcvt.s.d_b22-01.S",
  "rv64i_m/D/src/fcvt.s.d_b23-01.S",
  "rv64i_m/D/src/fcvt.s.d_b24-01.S",
  "rv64i_m/D/src/fcvt.s.d_b27-01.S",
  "rv64i_m/D/src/fcvt.s.d_b28-01.S",
  "rv64i_m/D/src/fcvt.s.d_b29-01.S",
  "rv64i_m/D/src/fcvt.w.d_b1-01.S",
  "rv64i_m/D/src/fcvt.w.d_b22-01.S",
  "rv64i_m/D/src/fcvt.w.d_b23-01.S",
  "rv64i_m/D/src/fcvt.w.d_b24-01.S",
  "rv64i_m/D/src/fcvt.w.d_b27-01.S",
  "rv64i_m/D/src/fcvt.w.d_b28-01.S",
  "rv64i_m/D/src/fcvt.w.d_b29-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b1-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b22-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b23-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b24-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b27-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b28-01.S",
  "rv64i_m/D/src/fcvt.wu.d_b29-01.S",
  "rv64i_m/D/src/feq.d_b1-01.S",
  "rv64i_m/D/src/feq.d_b19-01.S",
  "rv64i_m/D/src/fle.d_b1-01.S",
  "rv64i_m/D/src/fle.d_b19-01.S",
  "rv64i_m/D/src/flt.d_b1-01.S",
  "rv64i_m/D/src/flt.d_b19-01.S",
  "rv64i_m/D/src/fld-align-01.S",
  "rv64i_m/D/src/fsd-align-01.S",
  "rv64i_m/D/src/fmadd.d_b14-01.S",
  "rv64i_m/D/src/fmadd.d_b16-01.S",
  "rv64i_m/D/src/fmadd.d_b17-01.S",
  "rv64i_m/D/src/fmadd.d_b18-01.S",
  "rv64i_m/D/src/fmadd.d_b2-01.S",
  "rv64i_m/D/src/fmadd.d_b3-01.S",
  "rv64i_m/D/src/fmadd.d_b4-01.S",
  "rv64i_m/D/src/fmadd.d_b5-01.S",
  "rv64i_m/D/src/fmadd.d_b6-01.S",
  "rv64i_m/D/src/fmadd.d_b7-01.S",
  "rv64i_m/D/src/fmadd.d_b8-01.S",
  "rv64i_m/D/src/fmax.d_b1-01.S",
  "rv64i_m/D/src/fmax.d_b19-01.S",
  "rv64i_m/D/src/fmin.d_b1-01.S",
  "rv64i_m/D/src/fmin.d_b19-01.S",
  "rv64i_m/D/src/fmsub.d_b14-01.S",
  "rv64i_m/D/src/fmsub.d_b16-01.S",
  "rv64i_m/D/src/fmsub.d_b17-01.S",
  "rv64i_m/D/src/fmsub.d_b18-01.S",
  "rv64i_m/D/src/fmsub.d_b2-01.S",
  "rv64i_m/D/src/fmsub.d_b3-01.S",
  "rv64i_m/D/src/fmsub.d_b4-01.S",
  "rv64i_m/D/src/fmsub.d_b5-01.S",
  "rv64i_m/D/src/fmsub.d_b6-01.S",
  "rv64i_m/D/src/fmsub.d_b7-01.S",
  "rv64i_m/D/src/fmsub.d_b8-01.S",
  "rv64i_m/D/src/fmul.d_b1-01.S",
  "rv64i_m/D/src/fmul.d_b2-01.S",
  "rv64i_m/D/src/fmul.d_b3-01.S",
  "rv64i_m/D/src/fmul.d_b4-01.S",
  "rv64i_m/D/src/fmul.d_b5-01.S",
  "rv64i_m/D/src/fmul.d_b6-01.S",
  "rv64i_m/D/src/fmul.d_b7-01.S",
  "rv64i_m/D/src/fmul.d_b8-01.S",
  "rv64i_m/D/src/fmul.d_b9-01.S",
  "rv64i_m/D/src/fmv.d.x_b25-01.S",
  "rv64i_m/D/src/fmv.d.x_b26-01.S",
  "rv64i_m/D/src/fmv.x.d_b1-01.S",
  "rv64i_m/D/src/fmv.x.d_b22-01.S",
  "rv64i_m/D/src/fmv.x.d_b23-01.S",
  "rv64i_m/D/src/fmv.x.d_b24-01.S",
  "rv64i_m/D/src/fmv.x.d_b27-01.S",
  "rv64i_m/D/src/fmv.x.d_b28-01.S",
  "rv64i_m/D/src/fmv.x.d_b29-01.S",
  "rv64i_m/D/src/fnmadd.d_b14-01.S",
  "rv64i_m/D/src/fnmadd.d_b16-01.S",
  "rv64i_m/D/src/fnmadd.d_b17-01.S",
  "rv64i_m/D/src/fnmadd.d_b18-01.S",
  "rv64i_m/D/src/fnmadd.d_b2-01.S",
  "rv64i_m/D/src/fnmadd.d_b3-01.S",
  "rv64i_m/D/src/fnmadd.d_b4-01.S",
  "rv64i_m/D/src/fnmadd.d_b5-01.S",
  "rv64i_m/D/src/fnmadd.d_b6-01.S",
  "rv64i_m/D/src/fnmadd.d_b7-01.S",
  "rv64i_m/D/src/fnmadd.d_b8-01.S",
  "rv64i_m/D/src/fnmsub.d_b14-01.S",
  "rv64i_m/D/src/fnmsub.d_b16-01.S",
  "rv64i_m/D/src/fnmsub.d_b17-01.S",
  "rv64i_m/D/src/fnmsub.d_b18-01.S",
  "rv64i_m/D/src/fnmsub.d_b2-01.S",
  "rv64i_m/D/src/fnmsub.d_b3-01.S",
  "rv64i_m/D/src/fnmsub.d_b4-01.S",
  "rv64i_m/D/src/fnmsub.d_b5-01.S",
  "rv64i_m/D/src/fnmsub.d_b6-01.S",
  "rv64i_m/D/src/fnmsub.d_b7-01.S",
  "rv64i_m/D/src/fnmsub.d_b8-01.S",
  "rv64i_m/D/src/fsgnj.d_b1-01.S",
  "rv64i_m/D/src/fsgnjn.d_b1-01.S",
  "rv64i_m/D/src/fsgnjx.d_b1-01.S",
  "rv64i_m/D/src/fssub.d_b10-01.S",
  "rv64i_m/D/src/fssub.d_b1-01.S",
  "rv64i_m/D/src/fssub.d_b11-01.S",
  "rv64i_m/D/src/fssub.d_b12-01.S",
  "rv64i_m/D/src/fssub.d_b13-01.S",
  "rv64i_m/D/src/fssub.d_b2-01.S",
  "rv64i_m/D/src/fssub.d_b3-01.S",
  "rv64i_m/D/src/fssub.d_b4-01.S",
  "rv64i_m/D/src/fssub.d_b5-01.S",
  "rv64i_m/D/src/fssub.d_b7-01.S",
  "rv64i_m/D/src/fssub.d_b8-01.S"
};

string arch64zicboz[] = '{ // as of 12/17/23 presently cbo.zero is the only CMO instruction with riscv-arch-test support
  `RISCVARCHTEST,
  "rv64i_m/CMO/src/cbo.zero-01.S"
};

string arch32zicboz[] = '{ // as of 12/17/23 presently cbo.zero is the only CMO instruction with riscv-arch-test support
  `RISCVARCHTEST,
  "rv32i_m/CMO/src/cbo.zero-01.S"
};

string arch64zcb[] = '{
  `RISCVARCHTEST,
  "rv64i_m/C/src/clbu-01.S",
  "rv64i_m/C/src/clh-01.S",
  "rv64i_m/C/src/clhu-01.S",
  "rv64i_m/C/src/csb-01.S",
  "rv64i_m/C/src/csh-01.S",
  "rv64i_m/C/src/csext.b-01.S",
  "rv64i_m/C/src/csext.h-01.S",
  "rv64i_m/C/src/czext.b-01.S",
  "rv64i_m/C/src/czext.h-01.S",
  "rv64i_m/C/src/cmul-01.S",
  "rv64i_m/C/src/cnot-01.S",
  "rv64i_m/C/src/czext.w-01.S"
};

string arch32zcb[] = '{
  `RISCVARCHTEST,
  "rv32i_m/C/src/clbu-01.S",
  "rv32i_m/C/src/clh-01.S",
  "rv32i_m/C/src/clhu-01.S",
  "rv32i_m/C/src/csb-01.S",
  "rv32i_m/C/src/csh-01.S",
  "rv32i_m/C/src/csext.b-01.S",
  "rv32i_m/C/src/csext.h-01.S",
  "rv32i_m/C/src/czext.b-01.S",
  "rv32i_m/C/src/czext.h-01.S",
  "rv32i_m/C/src/cmul-01.S",
  "rv32i_m/C/src/cnot-01.S"
};

string arch64zba[] = '{
  `RISCVARCHTEST,
  "rv64i_m/B/src/slli.uw-01.S",
  "rv64i_m/B/src/add.uw-01.S",
  "rv64i_m/B/src/sh1add-01.S",
  "rv64i_m/B/src/sh2add-01.S",
  "rv64i_m/B/src/sh3add-01.S",
  "rv64i_m/B/src/sh1add.uw-01.S",
  "rv64i_m/B/src/sh2add.uw-01.S",
  "rv64i_m/B/src/sh3add.uw-01.S"
};

string arch64zbb[] = '{
  `RISCVARCHTEST,
  "rv64i_m/B/src/max-01.S",
  "rv64i_m/B/src/maxu-01.S",
  "rv64i_m/B/src/min-01.S",
  "rv64i_m/B/src/minu-01.S",
  "rv64i_m/B/src/orcb_64-01.S",
  "rv64i_m/B/src/rev8-01.S",
  "rv64i_m/B/src/andn-01.S",
  "rv64i_m/B/src/orn-01.S",
  "rv64i_m/B/src/xnor-01.S",
  "rv64i_m/B/src/zext.h_64-01.S",
  "rv64i_m/B/src/sext.b-01.S",
  "rv64i_m/B/src/sext.h-01.S",
  "rv64i_m/B/src/clz-01.S",
  "rv64i_m/B/src/clzw-01.S",
  "rv64i_m/B/src/cpop-01.S",
  "rv64i_m/B/src/cpopw-01.S",
  "rv64i_m/B/src/ctz-01.S",
  "rv64i_m/B/src/ctzw-01.S",
  "rv64i_m/B/src/rolw-01.S",
  "rv64i_m/B/src/ror-01.S",
  "rv64i_m/B/src/rori-01.S",
  "rv64i_m/B/src/roriw-01.S",
  "rv64i_m/B/src/rorw-01.S",
  "rv64i_m/B/src/rol-01.S"
};

string arch64zbc[] = '{
  `RISCVARCHTEST,
  "rv64i_m/B/src/clmul-01.S",
  "rv64i_m/B/src/clmulh-01.S",
  "rv64i_m/B/src/clmulr-01.S"
};

string arch64zbs[] = '{
  `RISCVARCHTEST,
  "rv64i_m/B/src/bclr-01.S",
  "rv64i_m/B/src/bclri-01.S",
  "rv64i_m/B/src/bext-01.S",
  "rv64i_m/B/src/bexti-01.S",
  "rv64i_m/B/src/binv-01.S",
  "rv64i_m/B/src/binvi-01.S",
  "rv64i_m/B/src/bset-01.S",
  "rv64i_m/B/src/bseti-01.S"
};

string arch64zbkc[] = '{
`RISCVARCHTEST,
"rv64i_m/B/src/clmul-01.S",
"rv64i_m/B/src/clmulh-01.S"
};

string arch64zbkx[] = '{
`RISCVARCHTEST,
"rv64i_m/K/src/xperm8-01.S",
"rv64i_m/K/src/xperm4-01.S"
};

string arch64zknd[] = '{
`RISCVARCHTEST,
"rv64i_m/K/src/aes64ds-01.S",
"rv64i_m/K/src/aes64dsm-01.S",
"rv64i_m/K/src/aes64im-01.S",
"rv64i_m/K/src/aes64ks1i-01.S",
"rv64i_m/K/src/aes64ks2-01.S"
};

string arch64zkne[] = '{
`RISCVARCHTEST,
"rv64i_m/K/src/aes64es-01.S",
"rv64i_m/K/src/aes64esm-01.S",
"rv64i_m/K/src/aes64ks1i-01.S",
"rv64i_m/K/src/aes64ks2-01.S"
};

string arch64zknh[] = '{
`RISCVARCHTEST,
"rv64i_m/K/src/sha256sig0-01.S",
"rv64i_m/K/src/sha256sig1-01.S",
"rv64i_m/K/src/sha256sum0-01.S",
"rv64i_m/K/src/sha256sum1-01.S",
"rv64i_m/K/src/sha512sig0-01.S",
"rv64i_m/K/src/sha512sig1-01.S",
"rv64i_m/K/src/sha512sum0-01.S",
"rv64i_m/K/src/sha512sum1-01.S"
};

string arch32priv[] = '{
  `RISCVARCHTEST,
  "rv32i_m/privilege/src/ebreak.S",
  "rv32i_m/privilege/src/ecall.S",
  "rv32i_m/privilege/src/misalign2-jalr-01.S",
  "rv32i_m/privilege/src/misalign-beq-01.S",
  "rv32i_m/privilege/src/misalign-bge-01.S",
  "rv32i_m/privilege/src/misalign-bgeu-01.S",
  "rv32i_m/privilege/src/misalign-blt-01.S",
  "rv32i_m/privilege/src/misalign-bltu-01.S",
  "rv32i_m/privilege/src/misalign-bne-01.S",
  "rv32i_m/privilege/src/misalign-jal-01.S",
  "rv32i_m/privilege/src/misalign-lh-01.S",
  "rv32i_m/privilege/src/misalign-lhu-01.S",
  "rv32i_m/privilege/src/misalign-lw-01.S",
  "rv32i_m/privilege/src/misalign-sh-01.S",
  "rv32i_m/privilege/src/misalign-sw-01.S"
};

string arch32m[] = '{
  `RISCVARCHTEST,
  "rv32i_m/M/src/div-01.S",
  "rv32i_m/M/src/divu-01.S",
  "rv32i_m/M/src/rem-01.S",
  "rv32i_m/M/src/remu-01.S",
  "rv32i_m/M/src/mul-01.S",
  "rv32i_m/M/src/mulh-01.S",
  "rv32i_m/M/src/mulhsu-01.S",
  "rv32i_m/M/src/mulhu-01.S"
};

string arch32f_fma[] = '{
  `RISCVARCHTEST,
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-001.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-002.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-003.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-004.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-005.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-006.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-007.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-008.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-009.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-010.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-011.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-012.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-013.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-014.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-015.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-016.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-017.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-018.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-019.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-020.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-021.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-022.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-023.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-024.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-025.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-026.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-027.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-028.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-029.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-030.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-031.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-032.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-033.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-034.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-035.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-036.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-037.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-038.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-039.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-040.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-041.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-042.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-043.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-044.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-045.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-046.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-047.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-048.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-049.S",
  // "rv32i_m/F/src/fmadd_b15/fmadd_b15-050.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-001.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-002.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-003.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-004.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-005.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-006.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-007.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-008.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-009.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-010.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-011.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-012.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-013.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-014.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-015.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-016.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-017.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-018.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-019.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-020.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-021.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-022.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-023.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-024.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-025.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-026.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-027.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-028.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-029.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-030.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-031.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-032.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-033.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-034.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-035.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-036.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-037.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-038.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-039.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-040.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-041.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-042.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-043.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-044.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-045.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-046.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-047.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-048.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-049.S",
  "rv32i_m/F/src/fmsub_b15/fmsub_b15-050.S"
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-001.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-002.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-003.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-004.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-005.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-006.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-007.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-008.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-009.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-010.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-011.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-012.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-013.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-014.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-015.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-016.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-017.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-018.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-019.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-020.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-021.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-022.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-023.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-024.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-025.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-026.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-027.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-028.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-029.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-030.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-031.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-032.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-033.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-034.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-035.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-036.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-037.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-038.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-039.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-040.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-041.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-042.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-043.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-044.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-045.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-046.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-047.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-048.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-049.S",
  // "rv32i_m/F/src/fnmadd_b15/fnmadd_b15-050.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-001.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-002.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-003.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-004.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-005.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-006.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-007.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-008.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-009.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-010.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-011.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-012.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-013.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-014.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-015.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-016.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-017.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-018.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-019.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-020.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-021.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-022.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-023.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-024.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-025.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-026.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-027.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-028.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-029.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-030.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-031.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-032.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-033.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-034.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-035.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-036.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-037.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-038.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-039.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-040.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-041.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-042.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-043.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-044.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-045.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-046.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-047.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-048.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-049.S",
  // "rv32i_m/F/src/fnmsub_b15/fnmsub_b15-050.S"
};

string arch32f_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv32i_m/F/src/fdiv_b20-01.S",
  "rv32i_m/F/src/fdiv_b1-01.S",
  "rv32i_m/F/src/fdiv_b2-01.S",
  "rv32i_m/F/src/fdiv_b21-01.S",
  "rv32i_m/F/src/fdiv_b3-01.S",
  "rv32i_m/F/src/fdiv_b4-01.S",
  "rv32i_m/F/src/fdiv_b5-01.S",
  "rv32i_m/F/src/fdiv_b6-01.S",
  "rv32i_m/F/src/fdiv_b7-01.S",
  "rv32i_m/F/src/fdiv_b8-01.S",
  "rv32i_m/F/src/fdiv_b9-01.S",
  "rv32i_m/F/src/fsqrt_b1-01.S",
  "rv32i_m/F/src/fsqrt_b20-01.S",
  "rv32i_m/F/src/fsqrt_b2-01.S",
  "rv32i_m/F/src/fsqrt_b3-01.S",
  "rv32i_m/F/src/fsqrt_b4-01.S",
  "rv32i_m/F/src/fsqrt_b5-01.S",
  "rv32i_m/F/src/fsqrt_b7-01.S",
  "rv32i_m/F/src/fsqrt_b8-01.S",
  "rv32i_m/F/src/fsqrt_b9-01.S"
};

string arch32f[] = '{
  `RISCVARCHTEST,
  "rv32i_m/F/src/fadd_b11-01.S",
  "rv32i_m/F/src/fadd_b10-01.S",
  "rv32i_m/F/src/fadd_b1-01.S",
  "rv32i_m/F/src/fadd_b11-01.S",
  "rv32i_m/F/src/fadd_b12-01.S",
  "rv32i_m/F/src/fadd_b13-01.S",
  "rv32i_m/F/src/fadd_b2-01.S",
  "rv32i_m/F/src/fadd_b3-01.S",
  "rv32i_m/F/src/fadd_b4-01.S",
  "rv32i_m/F/src/fadd_b5-01.S",
  "rv32i_m/F/src/fadd_b7-01.S",
  "rv32i_m/F/src/fadd_b8-01.S",
  "rv32i_m/F/src/fclass_b1-01.S",
  "rv32i_m/F/src/fcvt.s.w_b25-01.S",
  "rv32i_m/F/src/fcvt.s.w_b26-01.S",
  "rv32i_m/F/src/fcvt.s.wu_b25-01.S",
  "rv32i_m/F/src/fcvt.s.wu_b26-01.S",
  "rv32i_m/F/src/fcvt.w.s_b1-01.S",
  "rv32i_m/F/src/fcvt.w.s_b22-01.S",
  "rv32i_m/F/src/fcvt.w.s_b23-01.S",
  "rv32i_m/F/src/fcvt.w.s_b24-01.S",
  "rv32i_m/F/src/fcvt.w.s_b27-01.S",
  "rv32i_m/F/src/fcvt.w.s_b28-01.S",
  "rv32i_m/F/src/fcvt.w.s_b29-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b1-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b22-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b23-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b24-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b27-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b28-01.S",
  "rv32i_m/F/src/fcvt.wu.s_b29-01.S",
  "rv32i_m/F/src/feq_b1-01.S",
  "rv32i_m/F/src/feq_b19-01.S",
  "rv32i_m/F/src/fle_b1-01.S",
  "rv32i_m/F/src/fle_b19-01.S",
  "rv32i_m/F/src/flt_b1-01.S",
  "rv32i_m/F/src/flt_b19-01.S",
  "rv32i_m/F/src/flw-align-01.S",
  "rv32i_m/F/src/fmadd_b1-01.S",
  "rv32i_m/F/src/fmadd_b14-01.S",
  "rv32i_m/F/src/fmadd_b16-01.S",
  "rv32i_m/F/src/fmadd_b17-01.S",
  "rv32i_m/F/src/fmadd_b18-01.S",
  "rv32i_m/F/src/fmadd_b2-01.S",
  "rv32i_m/F/src/fmadd_b3-01.S",
  "rv32i_m/F/src/fmadd_b4-01.S",
  "rv32i_m/F/src/fmadd_b5-01.S",
  "rv32i_m/F/src/fmadd_b6-01.S",
  "rv32i_m/F/src/fmadd_b7-01.S",
  "rv32i_m/F/src/fmadd_b8-01.S",
  "rv32i_m/F/src/fmax_b1-01.S",
  "rv32i_m/F/src/fmax_b19-01.S",
  "rv32i_m/F/src/fmin_b1-01.S",
  "rv32i_m/F/src/fmin_b19-01.S",
  "rv32i_m/F/src/fmsub_b1-01.S",
  "rv32i_m/F/src/fmsub_b14-01.S",
  "rv32i_m/F/src/fmsub_b16-01.S",
  "rv32i_m/F/src/fmsub_b17-01.S",
  "rv32i_m/F/src/fmsub_b18-01.S",
  "rv32i_m/F/src/fmsub_b2-01.S",
  "rv32i_m/F/src/fmsub_b3-01.S",
  "rv32i_m/F/src/fmsub_b4-01.S",
  "rv32i_m/F/src/fmsub_b5-01.S",
  "rv32i_m/F/src/fmsub_b6-01.S",
  "rv32i_m/F/src/fmsub_b7-01.S",
  "rv32i_m/F/src/fmsub_b8-01.S",
  "rv32i_m/F/src/fmul_b1-01.S",
  "rv32i_m/F/src/fmul_b2-01.S",
  "rv32i_m/F/src/fmul_b3-01.S",
  "rv32i_m/F/src/fmul_b4-01.S",
  "rv32i_m/F/src/fmul_b5-01.S",
  "rv32i_m/F/src/fmul_b6-01.S",
  "rv32i_m/F/src/fmul_b7-01.S",
  "rv32i_m/F/src/fmul_b8-01.S",
  "rv32i_m/F/src/fmul_b9-01.S",
  "rv32i_m/F/src/fmv.w.x_b25-01.S",
  "rv32i_m/F/src/fmv.w.x_b26-01.S",
  "rv32i_m/F/src/fmv.x.w_b1-01.S",
  "rv32i_m/F/src/fmv.x.w_b22-01.S",
  "rv32i_m/F/src/fmv.x.w_b23-01.S",
  "rv32i_m/F/src/fmv.x.w_b24-01.S",
  "rv32i_m/F/src/fmv.x.w_b27-01.S",
  "rv32i_m/F/src/fmv.x.w_b28-01.S",
  "rv32i_m/F/src/fmv.x.w_b29-01.S",
  "rv32i_m/F/src/fnmadd_b1-01.S",
  "rv32i_m/F/src/fnmadd_b14-01.S",
  "rv32i_m/F/src/fnmadd_b16-01.S",
  "rv32i_m/F/src/fnmadd_b17-01.S",
  "rv32i_m/F/src/fnmadd_b18-01.S",
  "rv32i_m/F/src/fnmadd_b2-01.S",
  "rv32i_m/F/src/fnmadd_b3-01.S",
  "rv32i_m/F/src/fnmadd_b4-01.S",
  "rv32i_m/F/src/fnmadd_b5-01.S",
  "rv32i_m/F/src/fnmadd_b6-01.S",
  "rv32i_m/F/src/fnmadd_b7-01.S",
  "rv32i_m/F/src/fnmadd_b8-01.S",
  "rv32i_m/F/src/fnmsub_b1-01.S",
  "rv32i_m/F/src/fnmsub_b14-01.S",
  "rv32i_m/F/src/fnmsub_b16-01.S",
  "rv32i_m/F/src/fnmsub_b17-01.S",
  "rv32i_m/F/src/fnmsub_b18-01.S",
  "rv32i_m/F/src/fnmsub_b2-01.S",
  "rv32i_m/F/src/fnmsub_b3-01.S",
  "rv32i_m/F/src/fnmsub_b4-01.S",
  "rv32i_m/F/src/fnmsub_b5-01.S",
  "rv32i_m/F/src/fnmsub_b6-01.S",
  "rv32i_m/F/src/fnmsub_b7-01.S",
  "rv32i_m/F/src/fnmsub_b8-01.S",
  "rv32i_m/F/src/fsgnj_b1-01.S",
  "rv32i_m/F/src/fsgnjn_b1-01.S",
  "rv32i_m/F/src/fsgnjx_b1-01.S",
  "rv32i_m/F/src/fsub_b10-01.S",
  "rv32i_m/F/src/fsub_b1-01.S",
  "rv32i_m/F/src/fsub_b11-01.S",
  "rv32i_m/F/src/fsub_b12-01.S",
  "rv32i_m/F/src/fsub_b13-01.S",
  "rv32i_m/F/src/fsub_b2-01.S",
  "rv32i_m/F/src/fsub_b3-01.S",
  "rv32i_m/F/src/fsub_b4-01.S",
  "rv32i_m/F/src/fsub_b5-01.S",
  "rv32i_m/F/src/fsub_b7-01.S",
  "rv32i_m/F/src/fsub_b8-01.S",
  "rv32i_m/F/src/fsw-align-01.S"
};

string arch32zfh_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv32i_m/Zfh/src/fdiv_b20-01.S",
  "rv32i_m/Zfh/src/fdiv_b1-01.S",
  "rv32i_m/Zfh/src/fdiv_b2-01.S",
  "rv32i_m/Zfh/src/fdiv_b21-01.S",
  "rv32i_m/Zfh/src/fdiv_b3-01.S",
  "rv32i_m/Zfh/src/fdiv_b4-01.S",
  "rv32i_m/Zfh/src/fdiv_b5-01.S",
  "rv32i_m/Zfh/src/fdiv_b6-01.S",
  "rv32i_m/Zfh/src/fdiv_b7-01.S",
  "rv32i_m/Zfh/src/fdiv_b8-01.S",
  "rv32i_m/Zfh/src/fdiv_b9-01.S",
  "rv32i_m/Zfh/src/fsqrt_b1-01.S",
  "rv32i_m/Zfh/src/fsqrt_b20-01.S",
  "rv32i_m/Zfh/src/fsqrt_b2-01.S",
  "rv32i_m/Zfh/src/fsqrt_b3-01.S",
  "rv32i_m/Zfh/src/fsqrt_b4-01.S",
  "rv32i_m/Zfh/src/fsqrt_b5-01.S",
  "rv32i_m/Zfh/src/fsqrt_b7-01.S",
  "rv32i_m/Zfh/src/fsqrt_b8-01.S",
  "rv32i_m/Zfh/src/fsqrt_b9-01.S"
};

string arch32zfh[] = '{
  `RISCVARCHTEST,
  "rv32i_m/Zfh/src/fadd_b10-01.S",
  "rv32i_m/Zfh/src/fadd_b1-01.S",
  "rv32i_m/Zfh/src/fadd_b11-01.S",
  "rv32i_m/Zfh/src/fadd_b12-01.S",
  "rv32i_m/Zfh/src/fadd_b13-01.S",
  "rv32i_m/Zfh/src/fadd_b2-01.S",
  "rv32i_m/Zfh/src/fadd_b3-01.S",
  "rv32i_m/Zfh/src/fadd_b4-01.S",
  "rv32i_m/Zfh/src/fadd_b5-01.S",
  "rv32i_m/Zfh/src/fadd_b7-01.S",
  "rv32i_m/Zfh/src/fadd_b8-01.S",
  "rv32i_m/Zfh/src/fclass_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.h.s_b29-01.S",
  "rv32i_m/Zfh/src/fcvt.h.w_b25-01.S",
  "rv32i_m/Zfh/src/fcvt.h.w_b26-01.S",
  "rv32i_m/Zfh/src/fcvt.h.wu_b25-01.S",
  "rv32i_m/Zfh/src/fcvt.h.wu_b26-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.s.h_b29-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.w.h_b29-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.wu.h_b29-01.S",
  "rv32i_m/Zfh/src/feq_b1-01.S",
  "rv32i_m/Zfh/src/feq_b19-01.S",
  "rv32i_m/Zfh/src/fle_b1-01.S",
  "rv32i_m/Zfh/src/fle_b19-01.S",
  "rv32i_m/Zfh/src/flt_b1-01.S",
  "rv32i_m/Zfh/src/flt_b19-01.S",
  "rv32i_m/Zfh/src/flh-align-01.S",
  "rv32i_m/Zfh/src/fmax_b1-01.S",
  "rv32i_m/Zfh/src/fmax_b19-01.S",
  "rv32i_m/Zfh/src/fmin_b1-01.S",
  "rv32i_m/Zfh/src/fmin_b19-01.S",
  "rv32i_m/Zfh/src/fmul_b1-01.S",
  "rv32i_m/Zfh/src/fmul_b2-01.S",
  "rv32i_m/Zfh/src/fmul_b3-01.S",
  "rv32i_m/Zfh/src/fmul_b4-01.S",
  "rv32i_m/Zfh/src/fmul_b5-01.S",
  "rv32i_m/Zfh/src/fmul_b6-01.S",
  "rv32i_m/Zfh/src/fmul_b7-01.S",
  "rv32i_m/Zfh/src/fmul_b8-01.S",
  "rv32i_m/Zfh/src/fmul_b9-01.S",
  "rv32i_m/Zfh/src/fmv.h.x_b25-01.S",
  "rv32i_m/Zfh/src/fmv.h.x_b26-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b1-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b22-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b23-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b24-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b27-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b28-01.S",
  "rv32i_m/Zfh/src/fmv.x.h_b29-01.S",
  "rv32i_m/Zfh/src/fsgnj_b1-01.S",
  "rv32i_m/Zfh/src/fsgnjn_b1-01.S",
  "rv32i_m/Zfh/src/fsgnjx_b1-01.S",
  "rv32i_m/Zfh/src/fsub_b10-01.S",
  "rv32i_m/Zfh/src/fsub_b1-01.S",
  "rv32i_m/Zfh/src/fsub_b11-01.S",
  "rv32i_m/Zfh/src/fsub_b12-01.S",
  "rv32i_m/Zfh/src/fsub_b13-01.S",
  "rv32i_m/Zfh/src/fsub_b2-01.S",
  "rv32i_m/Zfh/src/fsub_b3-01.S",
  "rv32i_m/Zfh/src/fsub_b4-01.S",
  "rv32i_m/Zfh/src/fsub_b5-01.S",
  "rv32i_m/Zfh/src/fsub_b7-01.S",
  "rv32i_m/Zfh/src/fsub_b8-01.S",
  "rv32i_m/Zfh/src/fsh-align-01.S",
  "rv32i_m/Zfh/src/fmadd_b14-01.S",
  "rv32i_m/Zfh/src/fmadd_b16-01.S",
  "rv32i_m/Zfh/src/fmadd_b17-01.S",
  "rv32i_m/Zfh/src/fmadd_b18-01.S",
  "rv32i_m/Zfh/src/fmadd_b2-01.S",
  "rv32i_m/Zfh/src/fmadd_b3-01.S",
  "rv32i_m/Zfh/src/fmadd_b4-01.S",
  "rv32i_m/Zfh/src/fmadd_b5-01.S",
  "rv32i_m/Zfh/src/fmadd_b6-01.S",
  "rv32i_m/Zfh/src/fmadd_b7-01.S",
  "rv32i_m/Zfh/src/fmadd_b8-01.S",
  "rv32i_m/Zfh/src/fmsub_b14-01.S",
  "rv32i_m/Zfh/src/fmsub_b16-01.S",
  "rv32i_m/Zfh/src/fmsub_b17-01.S",
  "rv32i_m/Zfh/src/fmsub_b18-01.S",
  "rv32i_m/Zfh/src/fmsub_b2-01.S",
  "rv32i_m/Zfh/src/fmsub_b3-01.S",
  "rv32i_m/Zfh/src/fmsub_b4-01.S",
  "rv32i_m/Zfh/src/fmsub_b5-01.S",
  "rv32i_m/Zfh/src/fmsub_b6-01.S",
  "rv32i_m/Zfh/src/fmsub_b7-01.S",
  "rv32i_m/Zfh/src/fmsub_b8-01.S",
  "rv32i_m/Zfh/src/fnmadd_b14-01.S",
  "rv32i_m/Zfh/src/fnmadd_b16-01.S",
  "rv32i_m/Zfh/src/fnmadd_b17-01.S",
  "rv32i_m/Zfh/src/fnmadd_b18-01.S",
  "rv32i_m/Zfh/src/fnmadd_b2-01.S",
  "rv32i_m/Zfh/src/fnmadd_b3-01.S",
  "rv32i_m/Zfh/src/fnmadd_b4-01.S",
  "rv32i_m/Zfh/src/fnmadd_b5-01.S",
  "rv32i_m/Zfh/src/fnmadd_b6-01.S",
  "rv32i_m/Zfh/src/fnmadd_b7-01.S",
  "rv32i_m/Zfh/src/fnmadd_b8-01.S",
  "rv32i_m/Zfh/src/fnmsub_b14-01.S",
  "rv32i_m/Zfh/src/fnmsub_b16-01.S",
  "rv32i_m/Zfh/src/fnmsub_b17-01.S",
  "rv32i_m/Zfh/src/fnmsub_b18-01.S",
  "rv32i_m/Zfh/src/fnmsub_b2-01.S",
  "rv32i_m/Zfh/src/fnmsub_b3-01.S",
  "rv32i_m/Zfh/src/fnmsub_b4-01.S",
  "rv32i_m/Zfh/src/fnmsub_b5-01.S",
  "rv32i_m/Zfh/src/fnmsub_b6-01.S",
  "rv32i_m/Zfh/src/fnmsub_b7-01.S",
  "rv32i_m/Zfh/src/fnmsub_b8-01.S"
};

string arch32zfh_d[] = '{
  // `RISCVARCHTEST,
  "rv32i_m/Zfh/src/fcvt.d.h_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.d.h_b29-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b1-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b22-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b23-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b24-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b27-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b28-01.S",
  "rv32i_m/Zfh/src/fcvt.h.d_b29-01.S"
};

string arch32zfaf[] = '{
  `RISCVARCHTEST,
  "rv32i_m/F_Zfa/src/fround_b1-01.S",
  "rv32i_m/F_Zfa/src/froundnx_b1-01.S",
  "rv32i_m/F_Zfa/src/fleq_b1-01.S",
  "rv32i_m/F_Zfa/src/fleq_b19-01.S",
  "rv32i_m/F_Zfa/src/fli.s-01.S",
  "rv32i_m/F_Zfa/src/fltq_b1-01.S",
  "rv32i_m/F_Zfa/src/fltq_b19-01.S",
  "rv32i_m/D_Zfa/src/fltq_b1-01.S", // these D tests are more comprehensive and seem they should replace the F tests.  Applies to all F tests duplicated in D
  "rv32i_m/D_Zfa/src/fltq_b19-01.S",
  "rv32i_m/F_Zfa/src/fminm_b1-01.S",
  "rv32i_m/F_Zfa/src/fminm_b19-01.S",
  "rv32i_m/F_Zfa/src/fmaxm_b1-01.S",
  "rv32i_m/F_Zfa/src/fmaxm_b19-01.S"
};

string arch32zfad[] = '{
  `RISCVARCHTEST,
  "rv32i_m/D_Zfa/src/fround_b1-01.S",
  "rv32i_m/D_Zfa/src/froundnx_b1-01.S",
  "rv32i_m/D_Zfa/src/fround.d_b1-01.S",
  "rv32i_m/D_Zfa/src/froundnx.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b22-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b23-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b24-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b27-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b28-01.S",
  "rv32i_m/D_Zfa/src/fcvtmod.w.d_b29-01.S",
  "rv32i_m/D_Zfa/src/fleq_b1-01.S",
  "rv32i_m/D_Zfa/src/fleq_b19-01.S",
  "rv32i_m/D_Zfa/src/fleq.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fleq.d_b19-01.S",
  "rv32i_m/D_Zfa/src/fli.d-01.S",
  "rv32i_m/D_Zfa/src/fltq_b1-01.S",
  "rv32i_m/D_Zfa/src/fltq_b19-01.S",
  "rv32i_m/D_Zfa/src/fltq.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fltq.d_b19-01.S",
  "rv32i_m/D_Zfa/src/fminm_b1-01.S",
  "rv32i_m/D_Zfa/src/fminm_b19-01.S",
  "rv32i_m/D_Zfa/src/fminm.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fminm.d_b19-01.S",
  "rv32i_m/D_Zfa/src/fmaxm_b1-01.S",
  "rv32i_m/D_Zfa/src/fmaxm_b19-01.S",
  "rv32i_m/D_Zfa/src/fmaxm.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fmaxm.d_b19-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b1-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b22-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b23-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b24-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b27-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b28-01.S",
  "rv32i_m/D_Zfa/src/fmvh.x.d_b29-01.S"
};

string arch64zfaf[] = '{
  `RISCVARCHTEST,
  "rv64i_m/F_Zfa/src/fround_b1-01.S",
  "rv64i_m/F_Zfa/src/froundnx_b1-01.S",
  "rv64i_m/F_Zfa/src/fleq_b1-01.S",
  "rv64i_m/F_Zfa/src/fleq_b19-01.S",
  "rv64i_m/F_Zfa/src/fli.s-01.S",
  "rv64i_m/F_Zfa/src/fltq_b1-01.S",
  "rv64i_m/F_Zfa/src/fltq_b19-01.S",
  "rv64i_m/F_Zfa/src/fminm_b1-01.S",
  "rv64i_m/F_Zfa/src/fminm_b19-01.S",
  "rv64i_m/F_Zfa/src/fmaxm_b1-01.S",
  "rv64i_m/F_Zfa/src/fmaxm_b19-01.S"
};

string arch64zfad[] = '{
  `RISCVARCHTEST,
  "rv64i_m/D_Zfa/src/fround_b1-01.S",
  "rv64i_m/D_Zfa/src/froundnx_b1-01.S",
  "rv64i_m/D_Zfa/src/fround.d_b1-01.S",
  "rv64i_m/D_Zfa/src/froundnx.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b22-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b23-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b24-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b27-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b28-01.S",
  "rv64i_m/D_Zfa/src/fcvtmod.w.d_b29-01.S",
  "rv64i_m/D_Zfa/src/fleq_b1-01.S",
  "rv64i_m/D_Zfa/src/fleq_b19-01.S",
  "rv64i_m/D_Zfa/src/fleq.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fleq.d_b19-01.S",
  "rv64i_m/D_Zfa/src/fli.d-01.S",
  "rv64i_m/D_Zfa/src/fltq_b1-01.S",
  "rv64i_m/D_Zfa/src/fltq_b19-01.S",
  "rv64i_m/D_Zfa/src/fltq.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fltq.d_b19-01.S",
  "rv64i_m/D_Zfa/src/fminm_b1-01.S",
  "rv64i_m/D_Zfa/src/fminm_b19-01.S",
  "rv64i_m/D_Zfa/src/fminm.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fminm.d_b19-01.S",
  "rv64i_m/D_Zfa/src/fmaxm_b1-01.S",
  "rv64i_m/D_Zfa/src/fmaxm_b19-01.S",
  "rv64i_m/D_Zfa/src/fmaxm.d_b1-01.S",
  "rv64i_m/D_Zfa/src/fmaxm.d_b19-01.S"
};

string arch32d_fma[] = '{
  `RISCVARCHTEST,
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-001.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-002.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-003.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-004.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-005.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-006.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-007.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-008.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-009.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-010.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-011.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-012.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-013.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-014.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-015.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-016.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-017.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-018.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-019.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-020.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-021.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-022.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-023.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-024.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-025.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-026.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-027.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-028.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-029.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-030.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-031.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-032.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-033.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-034.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-035.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-036.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-037.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-038.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-039.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-040.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-041.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-042.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-043.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-044.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-045.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-046.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-047.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-048.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-049.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-050.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-051.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-052.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-053.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-054.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-055.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-056.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-057.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-058.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-059.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-060.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-061.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-062.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-063.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-064.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-065.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-066.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-067.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-068.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-069.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-070.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-071.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-072.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-073.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-074.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-075.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-076.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-077.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-078.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-079.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-080.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-081.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-082.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-083.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-084.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-085.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-086.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-087.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-088.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-089.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-090.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-091.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-092.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-093.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-094.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-095.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-096.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-097.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-098.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-099.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-100.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-101.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-102.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-103.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-104.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-105.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-106.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-107.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-108.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-109.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-110.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-111.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-112.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-113.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-114.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-115.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-116.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-117.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-118.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-119.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-120.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-121.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-122.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-123.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-124.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-125.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-126.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-127.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-128.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-129.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-130.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-131.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-132.S",
  // "rv32i_m/D/src/fmadd.d_b15/fmadd.d_b15-133.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-001.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-002.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-003.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-004.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-005.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-006.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-007.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-008.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-009.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-010.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-011.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-012.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-013.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-014.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-015.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-016.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-017.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-018.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-019.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-020.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-021.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-022.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-023.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-024.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-025.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-026.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-027.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-028.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-029.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-030.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-031.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-032.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-033.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-034.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-035.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-036.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-037.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-038.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-039.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-040.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-041.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-042.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-043.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-044.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-045.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-046.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-047.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-048.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-049.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-050.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-051.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-052.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-053.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-054.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-055.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-056.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-057.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-058.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-059.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-060.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-061.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-062.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-063.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-064.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-065.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-066.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-067.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-068.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-069.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-070.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-071.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-072.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-073.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-074.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-075.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-076.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-077.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-078.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-079.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-080.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-081.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-082.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-083.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-084.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-085.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-086.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-087.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-088.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-089.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-090.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-091.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-092.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-093.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-094.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-095.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-096.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-097.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-098.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-099.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-100.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-101.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-102.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-103.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-104.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-105.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-106.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-107.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-108.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-109.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-110.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-111.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-112.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-113.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-114.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-115.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-116.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-117.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-118.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-119.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-120.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-121.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-122.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-123.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-124.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-125.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-126.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-127.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-128.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-129.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-130.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-131.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-132.S",
  // "rv32i_m/D/src/fmsub.d_b15/fmsub.d_b15-133.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-001.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-002.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-003.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-004.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-005.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-006.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-007.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-008.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-009.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-010.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-011.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-012.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-013.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-014.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-015.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-016.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-017.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-018.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-019.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-020.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-021.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-022.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-023.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-024.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-025.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-026.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-027.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-028.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-029.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-030.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-031.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-032.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-033.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-034.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-035.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-036.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-037.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-038.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-039.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-040.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-041.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-042.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-043.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-044.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-045.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-046.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-047.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-048.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-049.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-050.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-051.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-052.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-053.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-054.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-055.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-056.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-057.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-058.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-059.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-060.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-061.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-062.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-063.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-064.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-065.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-066.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-067.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-068.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-069.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-070.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-071.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-072.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-073.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-074.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-075.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-076.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-077.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-078.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-079.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-080.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-081.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-082.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-083.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-084.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-085.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-086.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-087.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-088.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-089.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-090.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-091.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-092.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-093.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-094.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-095.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-096.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-097.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-098.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-099.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-100.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-101.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-102.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-103.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-104.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-105.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-106.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-107.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-108.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-109.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-110.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-111.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-112.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-113.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-114.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-115.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-116.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-117.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-118.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-119.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-120.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-121.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-122.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-123.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-124.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-125.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-126.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-127.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-128.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-129.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-130.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-131.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-132.S",
  // "rv32i_m/D/src/fnmadd.d_b15/fnmadd.d_b15-133.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-001.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-002.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-003.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-004.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-005.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-006.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-007.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-008.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-009.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-010.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-011.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-012.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-013.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-014.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-015.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-016.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-017.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-018.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-019.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-020.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-021.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-022.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-023.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-024.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-025.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-026.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-027.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-028.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-029.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-030.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-031.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-032.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-033.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-034.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-035.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-036.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-037.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-038.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-039.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-040.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-041.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-042.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-043.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-044.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-045.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-046.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-047.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-048.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-049.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-050.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-051.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-052.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-053.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-054.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-055.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-056.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-057.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-058.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-059.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-060.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-061.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-062.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-063.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-064.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-065.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-066.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-067.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-068.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-069.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-070.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-071.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-072.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-073.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-074.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-075.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-076.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-077.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-078.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-079.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-080.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-081.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-082.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-083.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-084.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-085.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-086.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-087.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-088.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-089.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-090.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-091.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-092.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-093.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-094.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-095.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-096.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-097.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-098.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-099.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-100.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-101.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-102.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-103.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-104.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-105.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-106.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-107.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-108.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-109.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-110.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-111.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-112.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-113.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-114.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-115.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-116.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-117.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-118.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-119.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-120.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-121.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-122.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-123.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-124.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-125.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-126.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-127.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-128.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-129.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-130.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-131.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-132.S",
  "rv32i_m/D/src/fnmsub.d_b15/fnmsub.d_b15-133.S"
};

string arch32zfh_fma[] = '{
  `RISCVARCHTEST,
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-001.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-002.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-003.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-004.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-005.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-006.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-007.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-008.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-009.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-010.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-011.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-012.S",
  "rv32i_m/Zfh/src/fmadd_b15/fmadd_b15-013.S",

  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-001.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-002.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-003.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-004.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-005.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-006.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-007.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-008.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-009.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-010.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-011.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-012.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-013.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-014.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-015.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-016.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-017.S",
  "rv32i_m/Zfh/src/fmadd_b1/fmadd_b1-018.S",

  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-001.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-002.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-003.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-004.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-005.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-006.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-007.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-008.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-009.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-010.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-011.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-012.S",
  "rv32i_m/Zfh/src/fmsub_b15/fmsub_b15-013.S",

  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-001.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-002.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-003.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-004.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-005.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-006.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-007.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-008.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-009.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-010.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-011.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-012.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-013.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-014.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-015.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-016.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-017.S",
  "rv32i_m/Zfh/src/fmsub_b1/fmsub_b1-018.S",

  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-001.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-002.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-003.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-004.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-005.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-006.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-007.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-008.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-009.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-010.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-011.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-012.S",
  "rv32i_m/Zfh/src/fnmadd_b15/fnmadd_b15-013.S",

  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-001.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-002.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-003.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-004.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-005.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-006.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-007.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-008.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-009.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-010.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-011.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-012.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-013.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-014.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-015.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-016.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-017.S",
  "rv32i_m/Zfh/src/fnmadd_b1/fnmadd_b1-018.S",

  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-001.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-002.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-003.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-004.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-005.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-006.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-007.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-008.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-009.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-010.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-011.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-012.S",
  "rv32i_m/Zfh/src/fnmsub_b15/fnmsub_b15-013.S",

  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-001.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-002.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-003.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-004.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-005.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-006.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-007.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-008.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-009.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-010.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-011.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-012.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-013.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-014.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-015.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-016.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-017.S",
  "rv32i_m/Zfh/src/fnmsub_b1/fnmsub_b1-018.S"
};

string arch32d_divsqrt[] = '{
  `RISCVARCHTEST,
  "rv32i_m/D/src/fdiv.d_b1-01.S",
  "rv32i_m/D/src/fdiv.d_b20-01.S",
  "rv32i_m/D/src/fdiv.d_b2-01.S",
  "rv32i_m/D/src/fdiv.d_b21-01.S",
  "rv32i_m/D/src/fdiv.d_b3-01.S",
  "rv32i_m/D/src/fdiv.d_b4-01.S",
  "rv32i_m/D/src/fdiv.d_b5-01.S",
  "rv32i_m/D/src/fdiv.d_b6-01.S",
  "rv32i_m/D/src/fdiv.d_b7-01.S",
  "rv32i_m/D/src/fdiv.d_b8-01.S",
  "rv32i_m/D/src/fdiv.d_b9-01.S",
  "rv32i_m/D/src/fsqrt.d_b1-01.S",
  "rv32i_m/D/src/fsqrt.d_b20-01.S",
  "rv32i_m/D/src/fsqrt.d_b2-01.S",
  "rv32i_m/D/src/fsqrt.d_b3-01.S",
  "rv32i_m/D/src/fsqrt.d_b4-01.S",
  "rv32i_m/D/src/fsqrt.d_b5-01.S",
  "rv32i_m/D/src/fsqrt.d_b7-01.S",
  "rv32i_m/D/src/fsqrt.d_b8-01.S",
  "rv32i_m/D/src/fsqrt.d_b9-01.S"
};

string arch32d[] = '{
  `RISCVARCHTEST,
  "rv32i_m/D/src/fadd.d_b10-01.S",
  "rv32i_m/D/src/fadd.d_b1-01.S",
  "rv32i_m/D/src/fadd.d_b11-01.S",
  "rv32i_m/D/src/fadd.d_b12-01.S",
  "rv32i_m/D/src/fadd.d_b13-01.S",
  "rv32i_m/D/src/fadd.d_b2-01.S",
  "rv32i_m/D/src/fadd.d_b3-01.S",
  "rv32i_m/D/src/fadd.d_b4-01.S",
  "rv32i_m/D/src/fadd.d_b5-01.S",
  "rv32i_m/D/src/fadd.d_b7-01.S",
  "rv32i_m/D/src/fadd.d_b8-01.S",
  "rv32i_m/D/src/fclass.d_b1-01.S",
  "rv32i_m/D/src/fcvt.d.s_b1-01.S",
  "rv32i_m/D/src/fcvt.d.s_b22-01.S",
  "rv32i_m/D/src/fcvt.d.s_b23-01.S",
  "rv32i_m/D/src/fcvt.d.s_b24-01.S",
  "rv32i_m/D/src/fcvt.d.s_b27-01.S",
  "rv32i_m/D/src/fcvt.d.s_b28-01.S",
  "rv32i_m/D/src/fcvt.d.s_b29-01.S",
  "rv32i_m/D/src/fcvt.d.w_b25-01.S",
  "rv32i_m/D/src/fcvt.d.w_b26-01.S",
  "rv32i_m/D/src/fcvt.d.wu_b25-01.S",
  "rv32i_m/D/src/fcvt.d.wu_b26-01.S",
  "rv32i_m/D/src/fcvt.s.d_b1-01.S",
  "rv32i_m/D/src/fcvt.s.d_b22-01.S",
  "rv32i_m/D/src/fcvt.s.d_b23-01.S",
  "rv32i_m/D/src/fcvt.s.d_b24-01.S",
  "rv32i_m/D/src/fcvt.s.d_b27-01.S",
  "rv32i_m/D/src/fcvt.s.d_b28-01.S",
  "rv32i_m/D/src/fcvt.s.d_b29-01.S",
  "rv32i_m/D/src/fcvt.w.d_b1-01.S",
  "rv32i_m/D/src/fcvt.w.d_b22-01.S",
  "rv32i_m/D/src/fcvt.w.d_b23-01.S",
  "rv32i_m/D/src/fcvt.w.d_b24-01.S",
  "rv32i_m/D/src/fcvt.w.d_b27-01.S",
  "rv32i_m/D/src/fcvt.w.d_b28-01.S",
  "rv32i_m/D/src/fcvt.w.d_b29-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b1-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b22-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b23-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b24-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b27-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b28-01.S",
  "rv32i_m/D/src/fcvt.wu.d_b29-01.S",
  "rv32i_m/D/src/feq.d_b1-01.S",
  "rv32i_m/D/src/feq.d_b19-01.S",
  "rv32i_m/D/src/fle.d_b1-01.S",
  "rv32i_m/D/src/fle.d_b19-01.S",
  "rv32i_m/D/src/flt.d_b1-01.S",
  "rv32i_m/D/src/flt.d_b19-01.S",
  "rv32i_m/D/src/fld-align-01.S",
  "rv32i_m/D/src/fsd-align-01.S",
  "rv32i_m/D/src/fmadd.d_b14-01.S",
  "rv32i_m/D/src/fmadd.d_b16-01.S",
  "rv32i_m/D/src/fmadd.d_b17-01.S",
  "rv32i_m/D/src/fmadd.d_b18-01.S",
  "rv32i_m/D/src/fmadd.d_b2-01.S",
  "rv32i_m/D/src/fmadd.d_b3-01.S",
  "rv32i_m/D/src/fmadd.d_b4-01.S",
  "rv32i_m/D/src/fmadd.d_b5-01.S",
  "rv32i_m/D/src/fmadd.d_b6-01.S",
  "rv32i_m/D/src/fmadd.d_b7-01.S",
  "rv32i_m/D/src/fmadd.d_b8-01.S",
  "rv32i_m/D/src/fmax.d_b1-01.S",
  "rv32i_m/D/src/fmax.d_b19-01.S",
  "rv32i_m/D/src/fmin.d_b1-01.S",
  "rv32i_m/D/src/fmin.d_b19-01.S",
  "rv32i_m/D/src/fmsub.d_b14-01.S",
  "rv32i_m/D/src/fmsub.d_b16-01.S",
  "rv32i_m/D/src/fmsub.d_b17-01.S",
  "rv32i_m/D/src/fmsub.d_b18-01.S",
  "rv32i_m/D/src/fmsub.d_b2-01.S",
  "rv32i_m/D/src/fmsub.d_b3-01.S",
  "rv32i_m/D/src/fmsub.d_b4-01.S",
  "rv32i_m/D/src/fmsub.d_b5-01.S",
  "rv32i_m/D/src/fmsub.d_b6-01.S",
  "rv32i_m/D/src/fmsub.d_b7-01.S",
  "rv32i_m/D/src/fmsub.d_b8-01.S",
  "rv32i_m/D/src/fmul.d_b1-01.S",
  "rv32i_m/D/src/fmul.d_b2-01.S",
  "rv32i_m/D/src/fmul.d_b3-01.S",
  "rv32i_m/D/src/fmul.d_b4-01.S",
  "rv32i_m/D/src/fmul.d_b5-01.S",
  "rv32i_m/D/src/fmul.d_b6-01.S",
  "rv32i_m/D/src/fmul.d_b7-01.S",
  "rv32i_m/D/src/fmul.d_b8-01.S",
  "rv32i_m/D/src/fmul.d_b9-01.S",
  "rv32i_m/D/src/fnmadd.d_b14-01.S",
  "rv32i_m/D/src/fnmadd.d_b16-01.S",
  "rv32i_m/D/src/fnmadd.d_b17-01.S",
  "rv32i_m/D/src/fnmadd.d_b18-01.S",
  "rv32i_m/D/src/fnmadd.d_b2-01.S",
  "rv32i_m/D/src/fnmadd.d_b3-01.S",
  "rv32i_m/D/src/fnmadd.d_b4-01.S",
  "rv32i_m/D/src/fnmadd.d_b5-01.S",
  "rv32i_m/D/src/fnmadd.d_b6-01.S",
  "rv32i_m/D/src/fnmadd.d_b7-01.S",
  "rv32i_m/D/src/fnmadd.d_b8-01.S",
  "rv32i_m/D/src/fnmsub.d_b14-01.S",
  "rv32i_m/D/src/fnmsub.d_b16-01.S",
  "rv32i_m/D/src/fnmsub.d_b17-01.S",
  "rv32i_m/D/src/fnmsub.d_b18-01.S",
  "rv32i_m/D/src/fnmsub.d_b2-01.S",
  "rv32i_m/D/src/fnmsub.d_b3-01.S",
  "rv32i_m/D/src/fnmsub.d_b4-01.S",
  "rv32i_m/D/src/fnmsub.d_b5-01.S",
  "rv32i_m/D/src/fnmsub.d_b6-01.S",
  "rv32i_m/D/src/fnmsub.d_b7-01.S",
  "rv32i_m/D/src/fnmsub.d_b8-01.S",
  "rv32i_m/D/src/fsgnj.d_b1-01.S",
  "rv32i_m/D/src/fsgnjn.d_b1-01.S",
  "rv32i_m/D/src/fsgnjx.d_b1-01.S",
  "rv32i_m/D/src/fssub.d_b10-01.S",
  "rv32i_m/D/src/fssub.d_b1-01.S",
  "rv32i_m/D/src/fssub.d_b11-01.S",
  "rv32i_m/D/src/fssub.d_b12-01.S",
  "rv32i_m/D/src/fssub.d_b13-01.S",
  "rv32i_m/D/src/fssub.d_b2-01.S",
  "rv32i_m/D/src/fssub.d_b3-01.S",
  "rv32i_m/D/src/fssub.d_b4-01.S",
  "rv32i_m/D/src/fssub.d_b5-01.S",
  "rv32i_m/D/src/fssub.d_b7-01.S",
  "rv32i_m/D/src/fssub.d_b8-01.S"
};


string arch32c[] = '{
  `RISCVARCHTEST,
  "rv32i_m/C/src/cadd-01.S",
  "rv32i_m/C/src/caddi-01.S",
  "rv32i_m/C/src/caddi16sp-01.S",
  "rv32i_m/C/src/caddi4spn-01.S",
  "rv32i_m/C/src/cand-01.S",
  "rv32i_m/C/src/candi-01.S",
  "rv32i_m/C/src/cbeqz-01.S",
  "rv32i_m/C/src/cbnez-01.S",
  "rv32i_m/C/src/cj-01.S",
  "rv32i_m/C/src/cjal-01.S",
  "rv32i_m/C/src/cjalr-01.S",
  "rv32i_m/C/src/cjr-01.S",
  "rv32i_m/C/src/cli-01.S",
  "rv32i_m/C/src/clui-01.S",
  "rv32i_m/C/src/clw-01.S",
  "rv32i_m/C/src/clwsp-01.S",
  "rv32i_m/C/src/cmv-01.S",
  "rv32i_m/C/src/cnop-01.S",
  "rv32i_m/C/src/cor-01.S",
  "rv32i_m/C/src/cslli-01.S",
  "rv32i_m/C/src/csrai-01.S",
  "rv32i_m/C/src/csrli-01.S",
  "rv32i_m/C/src/csub-01.S",
  "rv32i_m/C/src/csw-01.S",
  "rv32i_m/C/src/cswsp-01.S",
  "rv32i_m/C/src/cxor-01.S"
//  "rv32i_m/C/src/misalign1-cjalr-01.S", // no longer in repo
//"rv32i_m/C/src/misalign1-cjr-01.S"
};

string arch32cpriv[] = '{
  // `RISCVARCHTEST,
  "rv32i_m/C/src/cebreak-01.S"
};

string arch32zcf[] = '{
  // `RISCVARCHTEST,
  "rv32i_m/F_Zcf/src/c.flw-01.S",
  "rv32i_m/F_Zcf/src/c.flwsp-01.S",
  "rv32i_m/F_Zcf/src/c.fsw-01.S",
  "rv32i_m/F_Zcf/src/c.fswsp-01.S"
};

string arch32zcd[] = '{
  // `RISCVARCHTEST,
  "rv32i_m/D_Zcd/src/c.fld-01.S",
  "rv32i_m/D_Zcd/src/c.fldsp-01.S",
  "rv32i_m/D_Zcd/src/c.fsd-01.S",
  "rv32i_m/D_Zcd/src/c.fsdsp-01.S"
};

string arch32i[] = '{
  `RISCVARCHTEST,
  "rv32i_m/I/src/add-01.S",
  "rv32i_m/I/src/addi-01.S",
  "rv32i_m/I/src/and-01.S",
  "rv32i_m/I/src/andi-01.S",
  "rv32i_m/I/src/auipc-01.S",
  "rv32i_m/I/src/beq-01.S",
  "rv32i_m/I/src/bge-01.S",
  "rv32i_m/I/src/bgeu-01.S",
  "rv32i_m/I/src/blt-01.S",
  "rv32i_m/I/src/bltu-01.S",
  "rv32i_m/I/src/bne-01.S",
  "rv32i_m/I/src/fence-01.S",
  "rv32i_m/I/src/jal-01.S",
  "rv32i_m/I/src/jalr-01.S",
  "rv32i_m/I/src/lb-align-01.S",
  "rv32i_m/I/src/lbu-align-01.S",
  "rv32i_m/I/src/lh-align-01.S",
  "rv32i_m/I/src/lhu-align-01.S",
  "rv32i_m/I/src/lui-01.S",
  "rv32i_m/I/src/lw-align-01.S",
  "rv32i_m/I/src/or-01.S",
  "rv32i_m/I/src/ori-01.S",
  "rv32i_m/I/src/sb-align-01.S",
  "rv32i_m/I/src/sh-align-01.S",
  "rv32i_m/I/src/sll-01.S",
  "rv32i_m/I/src/slli-01.S",
  "rv32i_m/I/src/slt-01.S",
  "rv32i_m/I/src/slti-01.S",
  "rv32i_m/I/src/sltiu-01.S",
  "rv32i_m/I/src/sltu-01.S",
  "rv32i_m/I/src/sra-01.S",
  "rv32i_m/I/src/srai-01.S",
  "rv32i_m/I/src/srl-01.S",
  "rv32i_m/I/src/srli-01.S",
  "rv32i_m/I/src/sub-01.S",
  "rv32i_m/I/src/sw-align-01.S",
  "rv32i_m/I/src/xor-01.S",
  "rv32i_m/I/src/xori-01.S"
};

string arch32e[] = '{
  `RISCVARCHTEST,
  "rv32e_m/E/src/add-01.S",
  "rv32e_m/E/src/addi-01.S",
  "rv32e_m/E/src/and-01.S",
  "rv32e_m/E/src/andi-01.S",
  "rv32e_m/E/src/auipc-01.S",
  "rv32e_m/E/src/bge-01.S",
  "rv32e_m/E/src/bgeu-01.S",
  "rv32e_m/E/src/blt-01.S",
  "rv32e_m/E/src/bltu-01.S",
  "rv32e_m/E/src/bne-01.S",
  "rv32e_m/E/src/jal-01.S",
  "rv32e_m/E/src/jalr-01.S",
  "rv32e_m/E/src/lb-align-01.S",
  "rv32e_m/E/src/lbu-align-01.S",
  "rv32e_m/E/src/lh-align-01.S",
  "rv32e_m/E/src/lhu-align-01.S",
  "rv32e_m/E/src/lui-01.S",
  "rv32e_m/E/src/lw-align-01.S",
  "rv32e_m/E/src/or-01.S",
  "rv32e_m/E/src/ori-01.S",
  "rv32e_m/E/src/sb-align-01.S",
  "rv32e_m/E/src/sh-align-01.S",
  "rv32e_m/E/src/sll-01.S",
  "rv32e_m/E/src/slli-01.S",
  "rv32e_m/E/src/slt-01.S",
  "rv32e_m/E/src/slti-01.S",
  "rv32e_m/E/src/sltiu-01.S",
  "rv32e_m/E/src/sltu-01.S",
  "rv32e_m/E/src/sra-01.S",
  "rv32e_m/E/src/srai-01.S",
  "rv32e_m/E/src/srl-01.S",
  "rv32e_m/E/src/srli-01.S",
  "rv32e_m/E/src/sub-01.S",
  "rv32e_m/E/src/sw-align-01.S",
  "rv32e_m/E/src/xor-01.S",
  "rv32e_m/E/src/xori-01.S"
};

string wally64priv[] = '{
  `WALLYTEST,
  "rv64i_m/privilege/src/WALLY-minfo-01.S",
  "rv64i_m/privilege/src/WALLY-misaligned-access-01.S",
  "rv64i_m/privilege/src/WALLY-csr-permission-s-01.S",
  "rv64i_m/privilege/src/WALLY-cboz-01.S",
  "rv64i_m/privilege/src/WALLY-cbom-01.S",
  "rv64i_m/privilege/src/WALLY-csr-permission-u-01.S",
  "rv64i_m/privilege/src/WALLY-mie-01.S",
  "rv64i_m/privilege/src/WALLY-minfo-01.S",
  "rv64i_m/privilege/src/WALLY-misa-01.S",
  // "rv64i_m/privilege/src/WALLY-mmu-sv39-01.S",  // run this if SVADU_SUPPORTED = 0
  // "rv64i_m/privilege/src/WALLY-mmu-sv48-01.S",  // run this if SVADU_SUPPORTED = 0
  "rv64i_m/privilege/src/WALLY-mmu-sv39-svadu-svnapot-svpbmt-01.S",  // run this if SVADU_SUPPORTED = 1
  "rv64i_m/privilege/src/WALLY-mmu-sv48-svadu-01.S",  // run this if SVADU_SUPPORTED = 1
  "rv64i_m/privilege/src/WALLY-mtvec-01.S",
  "rv64i_m/privilege/src/WALLY-pma-01.S",
  "rv64i_m/privilege/src/WALLY-pmp-01.S",
  "rv64i_m/privilege/src/WALLY-sie-01.S",
  "rv64i_m/privilege/src/WALLY-status-mie-01.S",
  "rv64i_m/privilege/src/WALLY-status-sie-01.S",
  "rv64i_m/privilege/src/WALLY-status-tw-01.S",
  "rv64i_m/privilege/src/WALLY-status-tvm-01.S",
  "rv64i_m/privilege/src/WALLY-status-fp-enabled-01.S",
  "rv64i_m/privilege/src/WALLY-stvec-01.S",
  "rv64i_m/privilege/src/WALLY-trap-01.S",
  "rv64i_m/privilege/src/WALLY-trap-s-01.S",
  "rv64i_m/privilege/src/WALLY-trap-sret-01.S",
  "rv64i_m/privilege/src/WALLY-trap-u-01.S",
  "rv64i_m/privilege/src/WALLY-wfi-01.S",
  "rv64i_m/privilege/src/WALLY-endianness-01.S",
  "rv64i_m/privilege/src/WALLY-status-xlen-01.S",
  "rv64i_m/privilege/src/WALLY-satp-invalid-01.S"
};

string wally64periph[] = '{
  `WALLYTEST,
  "rv64i_m/privilege/src/WALLY-periph-01.S",
  "rv64i_m/privilege/src/WALLY-clint-01.S",
  "rv64i_m/privilege/src/WALLY-gpio-01.S",
  "rv64i_m/privilege/src/WALLY-plic-01.S",
  "rv64i_m/privilege/src/WALLY-plic-s-01.S",
  "rv64i_m/privilege/src/WALLY-uart-01.S",
  "rv64i_m/privilege/src/WALLY-spi-01.S"
};

string wally32priv[] = '{
  `WALLYTEST,
  "rv32i_m/privilege/src/WALLY-csr-permission-s-01.S",
  "rv32i_m/privilege/src/WALLY-csr-permission-u-01.S",
  // "rv32i_m/privilege/src/WALLY-cbom-01.S",
  "rv32i_m/privilege/src/WALLY-cboz-01.S",
  "rv32i_m/privilege/src/WALLY-mie-01.S",
  "rv32i_m/privilege/src/WALLY-minfo-01.S",
  "rv32i_m/privilege/src/WALLY-misa-01.S",
  // "rv32i_m/privilege/src/WALLY-mmu-sv32-01.S",    // run this if SVADU_SUPPORTED = 0
  "rv32i_m/privilege/src/WALLY-mmu-sv32-svadu-01.S", // run this if SVADU_SUPPORTED = 1
  "rv32i_m/privilege/src/WALLY-mtvec-01.S",
  "rv32i_m/privilege/src/WALLY-pma-01.S",
  "rv32i_m/privilege/src/WALLY-pmp-01.S",
  "rv32i_m/privilege/src/WALLY-sie-01.S",
  "rv32i_m/privilege/src/WALLY-status-mie-01.S",
  "rv32i_m/privilege/src/WALLY-status-sie-01.S",
  "rv32i_m/privilege/src/WALLY-status-tw-01.S",
  "rv32i_m/privilege/src/WALLY-status-tvm-01.S",
  "rv32i_m/privilege/src/WALLY-status-fp-enabled-01.S",
  "rv32i_m/privilege/src/WALLY-stvec-01.S",
  "rv32i_m/privilege/src/WALLY-trap-01.S",
  "rv32i_m/privilege/src/WALLY-trap-s-01.S",
  "rv32i_m/privilege/src/WALLY-trap-sret-01.S",
  "rv32i_m/privilege/src/WALLY-trap-u-01.S",
  "rv32i_m/privilege/src/WALLY-wfi-01.S",
  "rv32i_m/privilege/src/WALLY-endianness-01.S",
  "rv32i_m/privilege/src/WALLY-satp-invalid-01.S",
  // These peripherals are here instead of wally32periph because they don't work on rv32imc, which lacks a PMP register to configure
  "rv32i_m/privilege/src/WALLY-periph-s-01.S",
  "rv32i_m/privilege/src/WALLY-gpio-01.S",
  "rv32i_m/privilege/src/WALLY-clint-01.S",
  "rv32i_m/privilege/src/WALLY-uart-01.S",
  "rv32i_m/privilege/src/WALLY-plic-01.S",
  "rv32i_m/privilege/src/WALLY-plic-s-01.S",
  "rv32i_m/privilege/src/WALLY-spi-01.S"
};

string wally32periph[] = '{
  `WALLYTEST,
  "rv32i_m/privilege/src/WALLY-periph-01.S"
};

string fpga[] = '{
  `CUSTOM,
  "NULL"
};

string custom[] = '{
  `CUSTOM,
  "NULL"
};

string ahb64[] = '{
  `RISCVARCHTEST,
  "rv64i_m/F/src/fadd_b11-01.S"
};

string ahb32[] = '{
  `RISCVARCHTEST,
  "rv32i_m/F/src/fadd_b11-01.S"
};

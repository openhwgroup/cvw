// The following module make up the basic building blocks that
// are used by the cla64, cla_sub64, and cla52.

module INVBLOCK ( GIN, GOUT );
   
   input  GIN;
   output GOUT;
   
   assign GOUT =  ~ GIN;
   
endmodule // INVBLOCK


module XXOR1 ( A, B, GIN, SUM );
   
   input  A;
   input  B;
   input  GIN;
   output SUM;
   
   assign SUM = ( ~ (A ^ B)) ^ GIN;
   
endmodule // XXOR1


module BLOCK0 ( A, B, POUT, GOUT );
   
   input  A;
   input  B;
   output POUT;
   output GOUT;
   
   assign POUT =  ~ (A | B);
   assign GOUT =  ~ (A & B);
   
endmodule // BLOCK0


module BLOCK1 ( PIN1, PIN2, GIN1, GIN2, POUT, GOUT );
   
   input  PIN1;
   input  PIN2;
   input  GIN1;
   input  GIN2;
   output POUT;
   output GOUT;
   
   assign POUT =  ~ (PIN1 | PIN2);
   assign GOUT =  ~ (GIN2 & (PIN2 | GIN1));
   
endmodule // BLOCK1


module BLOCK2 ( PIN1, PIN2, GIN1, GIN2, POUT, GOUT );
   
   input  PIN1;
   input  PIN2;
   input  GIN1;
   input  GIN2;
   output POUT;
   output GOUT;
   
   assign POUT =  ~ (PIN1 & PIN2);
   assign GOUT =  ~ (GIN2 | (PIN2 & GIN1));
   
endmodule // BLOCK2


module BLOCK1A ( PIN2, GIN1, GIN2, GOUT );
   
   input  PIN2;
   input  GIN1;
   input  GIN2;
   output GOUT;
   
   assign GOUT =  ~ (GIN2 & (PIN2 | GIN1));
   
endmodule // BLOCK1A


module BLOCK2A ( PIN2, GIN1, GIN2, GOUT );
   
   input  PIN2;
   input  GIN1;
   input  GIN2;
   output GOUT;
   
   assign GOUT =  ~ (GIN2 | (PIN2 & GIN1));
   
endmodule
//***KEP all 0:63, 0:64 ect changed - changed due to lint warning
module PRESTAGE_64 ( A, B, CIN, POUT, GOUT );
   
   input  [63:0] A;
   input [63:0]  B;
   input 	 CIN;
   
   output [63:0] POUT;
   output [64:0] GOUT;
   
   BLOCK0 U10 (A[0] , B[0] , POUT[0] , GOUT[1] );
   BLOCK0 U11 (A[1] , B[1] , POUT[1] , GOUT[2] );
   BLOCK0 U12 (A[2] , B[2] , POUT[2] , GOUT[3] );
   BLOCK0 U13 (A[3] , B[3] , POUT[3] , GOUT[4] );
   BLOCK0 U14 (A[4] , B[4] , POUT[4] , GOUT[5] );
   BLOCK0 U15 (A[5] , B[5] , POUT[5] , GOUT[6] );
   BLOCK0 U16 (A[6] , B[6] , POUT[6] , GOUT[7] );
   BLOCK0 U17 (A[7] , B[7] , POUT[7] , GOUT[8] );
   BLOCK0 U18 (A[8] , B[8] , POUT[8] , GOUT[9] );
   BLOCK0 U19 (A[9] , B[9] , POUT[9] , GOUT[10] );
   BLOCK0 U110 (A[10] , B[10] , POUT[10] , GOUT[11] );
   BLOCK0 U111 (A[11] , B[11] , POUT[11] , GOUT[12] );
   BLOCK0 U112 (A[12] , B[12] , POUT[12] , GOUT[13] );
   BLOCK0 U113 (A[13] , B[13] , POUT[13] , GOUT[14] );
   BLOCK0 U114 (A[14] , B[14] , POUT[14] , GOUT[15] );
   BLOCK0 U115 (A[15] , B[15] , POUT[15] , GOUT[16] );
   BLOCK0 U116 (A[16] , B[16] , POUT[16] , GOUT[17] );
   BLOCK0 U117 (A[17] , B[17] , POUT[17] , GOUT[18] );
   BLOCK0 U118 (A[18] , B[18] , POUT[18] , GOUT[19] );
   BLOCK0 U119 (A[19] , B[19] , POUT[19] , GOUT[20] );
   BLOCK0 U120 (A[20] , B[20] , POUT[20] , GOUT[21] );
   BLOCK0 U121 (A[21] , B[21] , POUT[21] , GOUT[22] );
   BLOCK0 U122 (A[22] , B[22] , POUT[22] , GOUT[23] );
   BLOCK0 U123 (A[23] , B[23] , POUT[23] , GOUT[24] );
   BLOCK0 U124 (A[24] , B[24] , POUT[24] , GOUT[25] );
   BLOCK0 U125 (A[25] , B[25] , POUT[25] , GOUT[26] );
   BLOCK0 U126 (A[26] , B[26] , POUT[26] , GOUT[27] );
   BLOCK0 U127 (A[27] , B[27] , POUT[27] , GOUT[28] );
   BLOCK0 U128 (A[28] , B[28] , POUT[28] , GOUT[29] );
   BLOCK0 U129 (A[29] , B[29] , POUT[29] , GOUT[30] );
   BLOCK0 U130 (A[30] , B[30] , POUT[30] , GOUT[31] );
   BLOCK0 U131 (A[31] , B[31] , POUT[31] , GOUT[32] );
   BLOCK0 U132 (A[32] , B[32] , POUT[32] , GOUT[33] );
   BLOCK0 U133 (A[33] , B[33] , POUT[33] , GOUT[34] );
   BLOCK0 U134 (A[34] , B[34] , POUT[34] , GOUT[35] );
   BLOCK0 U135 (A[35] , B[35] , POUT[35] , GOUT[36] );
   BLOCK0 U136 (A[36] , B[36] , POUT[36] , GOUT[37] );
   BLOCK0 U137 (A[37] , B[37] , POUT[37] , GOUT[38] );
   BLOCK0 U138 (A[38] , B[38] , POUT[38] , GOUT[39] );
   BLOCK0 U139 (A[39] , B[39] , POUT[39] , GOUT[40] );
   BLOCK0 U140 (A[40] , B[40] , POUT[40] , GOUT[41] );
   BLOCK0 U141 (A[41] , B[41] , POUT[41] , GOUT[42] );
   BLOCK0 U142 (A[42] , B[42] , POUT[42] , GOUT[43] );
   BLOCK0 U143 (A[43] , B[43] , POUT[43] , GOUT[44] );
   BLOCK0 U144 (A[44] , B[44] , POUT[44] , GOUT[45] );
   BLOCK0 U145 (A[45] , B[45] , POUT[45] , GOUT[46] );
   BLOCK0 U146 (A[46] , B[46] , POUT[46] , GOUT[47] );
   BLOCK0 U147 (A[47] , B[47] , POUT[47] , GOUT[48] );
   BLOCK0 U148 (A[48] , B[48] , POUT[48] , GOUT[49] );
   BLOCK0 U149 (A[49] , B[49] , POUT[49] , GOUT[50] );
   BLOCK0 U150 (A[50] , B[50] , POUT[50] , GOUT[51] );
   BLOCK0 U151 (A[51] , B[51] , POUT[51] , GOUT[52] );
   BLOCK0 U152 (A[52] , B[52] , POUT[52] , GOUT[53] );
   BLOCK0 U153 (A[53] , B[53] , POUT[53] , GOUT[54] );
   BLOCK0 U154 (A[54] , B[54] , POUT[54] , GOUT[55] );
   BLOCK0 U155 (A[55] , B[55] , POUT[55] , GOUT[56] );
   BLOCK0 U156 (A[56] , B[56] , POUT[56] , GOUT[57] );
   BLOCK0 U157 (A[57] , B[57] , POUT[57] , GOUT[58] );
   BLOCK0 U158 (A[58] , B[58] , POUT[58] , GOUT[59] );
   BLOCK0 U159 (A[59] , B[59] , POUT[59] , GOUT[60] );
   BLOCK0 U160 (A[60] , B[60] , POUT[60] , GOUT[61] );
   BLOCK0 U161 (A[61] , B[61] , POUT[61] , GOUT[62] );
   BLOCK0 U162 (A[62] , B[62] , POUT[62] , GOUT[63] );
   BLOCK0 U163 (A[63] , B[63] , POUT[63] , GOUT[64] );
   INVBLOCK U2 (CIN , GOUT[0] );
   
endmodule // PRESTAGE_64


module DBLC_0_64 ( PIN, GIN, POUT, GOUT );
   
   input  [63:0] PIN;
   input [64:0]  GIN;
   
   output [62:0] POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   BLOCK1A U21 (PIN[0] , GIN[0] , GIN[1] , GOUT[1] );
   BLOCK1 U32 (PIN[0] , PIN[1] , GIN[1] , GIN[2] , POUT[0] , GOUT[2] );
   BLOCK1 U33 (PIN[1] , PIN[2] , GIN[2] , GIN[3] , POUT[1] , GOUT[3] );
   BLOCK1 U34 (PIN[2] , PIN[3] , GIN[3] , GIN[4] , POUT[2] , GOUT[4] );
   BLOCK1 U35 (PIN[3] , PIN[4] , GIN[4] , GIN[5] , POUT[3] , GOUT[5] );
   BLOCK1 U36 (PIN[4] , PIN[5] , GIN[5] , GIN[6] , POUT[4] , GOUT[6] );
   BLOCK1 U37 (PIN[5] , PIN[6] , GIN[6] , GIN[7] , POUT[5] , GOUT[7] );
   BLOCK1 U38 (PIN[6] , PIN[7] , GIN[7] , GIN[8] , POUT[6] , GOUT[8] );
   BLOCK1 U39 (PIN[7] , PIN[8] , GIN[8] , GIN[9] , POUT[7] , GOUT[9] );
   BLOCK1 U310 (PIN[8] , PIN[9] , GIN[9] , GIN[10] , POUT[8] , GOUT[10] );
   BLOCK1 U311 (PIN[9] , PIN[10] , GIN[10] , GIN[11] , POUT[9] , GOUT[11] );
   BLOCK1 U312 (PIN[10] , PIN[11] , GIN[11] , GIN[12] , POUT[10] , GOUT[12] );
   BLOCK1 U313 (PIN[11] , PIN[12] , GIN[12] , GIN[13] , POUT[11] , GOUT[13] );
   BLOCK1 U314 (PIN[12] , PIN[13] , GIN[13] , GIN[14] , POUT[12] , GOUT[14] );
   BLOCK1 U315 (PIN[13] , PIN[14] , GIN[14] , GIN[15] , POUT[13] , GOUT[15] );
   BLOCK1 U316 (PIN[14] , PIN[15] , GIN[15] , GIN[16] , POUT[14] , GOUT[16] );
   BLOCK1 U317 (PIN[15] , PIN[16] , GIN[16] , GIN[17] , POUT[15] , GOUT[17] );
   BLOCK1 U318 (PIN[16] , PIN[17] , GIN[17] , GIN[18] , POUT[16] , GOUT[18] );
   BLOCK1 U319 (PIN[17] , PIN[18] , GIN[18] , GIN[19] , POUT[17] , GOUT[19] );
   BLOCK1 U320 (PIN[18] , PIN[19] , GIN[19] , GIN[20] , POUT[18] , GOUT[20] );
   BLOCK1 U321 (PIN[19] , PIN[20] , GIN[20] , GIN[21] , POUT[19] , GOUT[21] );
   BLOCK1 U322 (PIN[20] , PIN[21] , GIN[21] , GIN[22] , POUT[20] , GOUT[22] );
   BLOCK1 U323 (PIN[21] , PIN[22] , GIN[22] , GIN[23] , POUT[21] , GOUT[23] );
   BLOCK1 U324 (PIN[22] , PIN[23] , GIN[23] , GIN[24] , POUT[22] , GOUT[24] );
   BLOCK1 U325 (PIN[23] , PIN[24] , GIN[24] , GIN[25] , POUT[23] , GOUT[25] );
   BLOCK1 U326 (PIN[24] , PIN[25] , GIN[25] , GIN[26] , POUT[24] , GOUT[26] );
   BLOCK1 U327 (PIN[25] , PIN[26] , GIN[26] , GIN[27] , POUT[25] , GOUT[27] );
   BLOCK1 U328 (PIN[26] , PIN[27] , GIN[27] , GIN[28] , POUT[26] , GOUT[28] );
   BLOCK1 U329 (PIN[27] , PIN[28] , GIN[28] , GIN[29] , POUT[27] , GOUT[29] );
   BLOCK1 U330 (PIN[28] , PIN[29] , GIN[29] , GIN[30] , POUT[28] , GOUT[30] );
   BLOCK1 U331 (PIN[29] , PIN[30] , GIN[30] , GIN[31] , POUT[29] , GOUT[31] );
   BLOCK1 U332 (PIN[30] , PIN[31] , GIN[31] , GIN[32] , POUT[30] , GOUT[32] );
   BLOCK1 U333 (PIN[31] , PIN[32] , GIN[32] , GIN[33] , POUT[31] , GOUT[33] );
   BLOCK1 U334 (PIN[32] , PIN[33] , GIN[33] , GIN[34] , POUT[32] , GOUT[34] );
   BLOCK1 U335 (PIN[33] , PIN[34] , GIN[34] , GIN[35] , POUT[33] , GOUT[35] );
   BLOCK1 U336 (PIN[34] , PIN[35] , GIN[35] , GIN[36] , POUT[34] , GOUT[36] );
   BLOCK1 U337 (PIN[35] , PIN[36] , GIN[36] , GIN[37] , POUT[35] , GOUT[37] );
   BLOCK1 U338 (PIN[36] , PIN[37] , GIN[37] , GIN[38] , POUT[36] , GOUT[38] );
   BLOCK1 U339 (PIN[37] , PIN[38] , GIN[38] , GIN[39] , POUT[37] , GOUT[39] );
   BLOCK1 U340 (PIN[38] , PIN[39] , GIN[39] , GIN[40] , POUT[38] , GOUT[40] );
   BLOCK1 U341 (PIN[39] , PIN[40] , GIN[40] , GIN[41] , POUT[39] , GOUT[41] );
   BLOCK1 U342 (PIN[40] , PIN[41] , GIN[41] , GIN[42] , POUT[40] , GOUT[42] );
   BLOCK1 U343 (PIN[41] , PIN[42] , GIN[42] , GIN[43] , POUT[41] , GOUT[43] );
   BLOCK1 U344 (PIN[42] , PIN[43] , GIN[43] , GIN[44] , POUT[42] , GOUT[44] );
   BLOCK1 U345 (PIN[43] , PIN[44] , GIN[44] , GIN[45] , POUT[43] , GOUT[45] );
   BLOCK1 U346 (PIN[44] , PIN[45] , GIN[45] , GIN[46] , POUT[44] , GOUT[46] );
   BLOCK1 U347 (PIN[45] , PIN[46] , GIN[46] , GIN[47] , POUT[45] , GOUT[47] );
   BLOCK1 U348 (PIN[46] , PIN[47] , GIN[47] , GIN[48] , POUT[46] , GOUT[48] );
   BLOCK1 U349 (PIN[47] , PIN[48] , GIN[48] , GIN[49] , POUT[47] , GOUT[49] );
   BLOCK1 U350 (PIN[48] , PIN[49] , GIN[49] , GIN[50] , POUT[48] , GOUT[50] );
   BLOCK1 U351 (PIN[49] , PIN[50] , GIN[50] , GIN[51] , POUT[49] , GOUT[51] );
   BLOCK1 U352 (PIN[50] , PIN[51] , GIN[51] , GIN[52] , POUT[50] , GOUT[52] );
   BLOCK1 U353 (PIN[51] , PIN[52] , GIN[52] , GIN[53] , POUT[51] , GOUT[53] );
   BLOCK1 U354 (PIN[52] , PIN[53] , GIN[53] , GIN[54] , POUT[52] , GOUT[54] );
   BLOCK1 U355 (PIN[53] , PIN[54] , GIN[54] , GIN[55] , POUT[53] , GOUT[55] );
   BLOCK1 U356 (PIN[54] , PIN[55] , GIN[55] , GIN[56] , POUT[54] , GOUT[56] );
   BLOCK1 U357 (PIN[55] , PIN[56] , GIN[56] , GIN[57] , POUT[55] , GOUT[57] );
   BLOCK1 U358 (PIN[56] , PIN[57] , GIN[57] , GIN[58] , POUT[56] , GOUT[58] );
   BLOCK1 U359 (PIN[57] , PIN[58] , GIN[58] , GIN[59] , POUT[57] , GOUT[59] );
   BLOCK1 U360 (PIN[58] , PIN[59] , GIN[59] , GIN[60] , POUT[58] , GOUT[60] );
   BLOCK1 U361 (PIN[59] , PIN[60] , GIN[60] , GIN[61] , POUT[59] , GOUT[61] );
   BLOCK1 U362 (PIN[60] , PIN[61] , GIN[61] , GIN[62] , POUT[60] , GOUT[62] );
   BLOCK1 U363 (PIN[61] , PIN[62] , GIN[62] , GIN[63] , POUT[61] , GOUT[63] );
   BLOCK1 U364 (PIN[62] , PIN[63] , GIN[63] , GIN[64] , POUT[62] , GOUT[64] );
   
endmodule // DBLC_0_64


module DBLC_1_64 ( PIN, GIN, POUT, GOUT );
   
   input  [62:0] PIN;
   input [64:0]  GIN;
   
   output [60:0] POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   INVBLOCK U11 (GIN[1] , GOUT[1] );
   BLOCK2A U22 (PIN[0] , GIN[0] , GIN[2] , GOUT[2] );
   BLOCK2A U23 (PIN[1] , GIN[1] , GIN[3] , GOUT[3] );
   BLOCK2 U34 (PIN[0] , PIN[2] , GIN[2] , GIN[4] , POUT[0] , GOUT[4] );
   BLOCK2 U35 (PIN[1] , PIN[3] , GIN[3] , GIN[5] , POUT[1] , GOUT[5] );
   BLOCK2 U36 (PIN[2] , PIN[4] , GIN[4] , GIN[6] , POUT[2] , GOUT[6] );
   BLOCK2 U37 (PIN[3] , PIN[5] , GIN[5] , GIN[7] , POUT[3] , GOUT[7] );
   BLOCK2 U38 (PIN[4] , PIN[6] , GIN[6] , GIN[8] , POUT[4] , GOUT[8] );
   BLOCK2 U39 (PIN[5] , PIN[7] , GIN[7] , GIN[9] , POUT[5] , GOUT[9] );
   BLOCK2 U310 (PIN[6] , PIN[8] , GIN[8] , GIN[10] , POUT[6] , GOUT[10] );
   BLOCK2 U311 (PIN[7] , PIN[9] , GIN[9] , GIN[11] , POUT[7] , GOUT[11] );
   BLOCK2 U312 (PIN[8] , PIN[10] , GIN[10] , GIN[12] , POUT[8] , GOUT[12] );
   BLOCK2 U313 (PIN[9] , PIN[11] , GIN[11] , GIN[13] , POUT[9] , GOUT[13] );
   BLOCK2 U314 (PIN[10] , PIN[12] , GIN[12] , GIN[14] , POUT[10] , GOUT[14] );
   BLOCK2 U315 (PIN[11] , PIN[13] , GIN[13] , GIN[15] , POUT[11] , GOUT[15] );
   BLOCK2 U316 (PIN[12] , PIN[14] , GIN[14] , GIN[16] , POUT[12] , GOUT[16] );
   BLOCK2 U317 (PIN[13] , PIN[15] , GIN[15] , GIN[17] , POUT[13] , GOUT[17] );
   BLOCK2 U318 (PIN[14] , PIN[16] , GIN[16] , GIN[18] , POUT[14] , GOUT[18] );
   BLOCK2 U319 (PIN[15] , PIN[17] , GIN[17] , GIN[19] , POUT[15] , GOUT[19] );
   BLOCK2 U320 (PIN[16] , PIN[18] , GIN[18] , GIN[20] , POUT[16] , GOUT[20] );
   BLOCK2 U321 (PIN[17] , PIN[19] , GIN[19] , GIN[21] , POUT[17] , GOUT[21] );
   BLOCK2 U322 (PIN[18] , PIN[20] , GIN[20] , GIN[22] , POUT[18] , GOUT[22] );
   BLOCK2 U323 (PIN[19] , PIN[21] , GIN[21] , GIN[23] , POUT[19] , GOUT[23] );
   BLOCK2 U324 (PIN[20] , PIN[22] , GIN[22] , GIN[24] , POUT[20] , GOUT[24] );
   BLOCK2 U325 (PIN[21] , PIN[23] , GIN[23] , GIN[25] , POUT[21] , GOUT[25] );
   BLOCK2 U326 (PIN[22] , PIN[24] , GIN[24] , GIN[26] , POUT[22] , GOUT[26] );
   BLOCK2 U327 (PIN[23] , PIN[25] , GIN[25] , GIN[27] , POUT[23] , GOUT[27] );
   BLOCK2 U328 (PIN[24] , PIN[26] , GIN[26] , GIN[28] , POUT[24] , GOUT[28] );
   BLOCK2 U329 (PIN[25] , PIN[27] , GIN[27] , GIN[29] , POUT[25] , GOUT[29] );
   BLOCK2 U330 (PIN[26] , PIN[28] , GIN[28] , GIN[30] , POUT[26] , GOUT[30] );
   BLOCK2 U331 (PIN[27] , PIN[29] , GIN[29] , GIN[31] , POUT[27] , GOUT[31] );
   BLOCK2 U332 (PIN[28] , PIN[30] , GIN[30] , GIN[32] , POUT[28] , GOUT[32] );
   BLOCK2 U333 (PIN[29] , PIN[31] , GIN[31] , GIN[33] , POUT[29] , GOUT[33] );
   BLOCK2 U334 (PIN[30] , PIN[32] , GIN[32] , GIN[34] , POUT[30] , GOUT[34] );
   BLOCK2 U335 (PIN[31] , PIN[33] , GIN[33] , GIN[35] , POUT[31] , GOUT[35] );
   BLOCK2 U336 (PIN[32] , PIN[34] , GIN[34] , GIN[36] , POUT[32] , GOUT[36] );
   BLOCK2 U337 (PIN[33] , PIN[35] , GIN[35] , GIN[37] , POUT[33] , GOUT[37] );
   BLOCK2 U338 (PIN[34] , PIN[36] , GIN[36] , GIN[38] , POUT[34] , GOUT[38] );
   BLOCK2 U339 (PIN[35] , PIN[37] , GIN[37] , GIN[39] , POUT[35] , GOUT[39] );
   BLOCK2 U340 (PIN[36] , PIN[38] , GIN[38] , GIN[40] , POUT[36] , GOUT[40] );
   BLOCK2 U341 (PIN[37] , PIN[39] , GIN[39] , GIN[41] , POUT[37] , GOUT[41] );
   BLOCK2 U342 (PIN[38] , PIN[40] , GIN[40] , GIN[42] , POUT[38] , GOUT[42] );
   BLOCK2 U343 (PIN[39] , PIN[41] , GIN[41] , GIN[43] , POUT[39] , GOUT[43] );
   BLOCK2 U344 (PIN[40] , PIN[42] , GIN[42] , GIN[44] , POUT[40] , GOUT[44] );
   BLOCK2 U345 (PIN[41] , PIN[43] , GIN[43] , GIN[45] , POUT[41] , GOUT[45] );
   BLOCK2 U346 (PIN[42] , PIN[44] , GIN[44] , GIN[46] , POUT[42] , GOUT[46] );
   BLOCK2 U347 (PIN[43] , PIN[45] , GIN[45] , GIN[47] , POUT[43] , GOUT[47] );
   BLOCK2 U348 (PIN[44] , PIN[46] , GIN[46] , GIN[48] , POUT[44] , GOUT[48] );
   BLOCK2 U349 (PIN[45] , PIN[47] , GIN[47] , GIN[49] , POUT[45] , GOUT[49] );
   BLOCK2 U350 (PIN[46] , PIN[48] , GIN[48] , GIN[50] , POUT[46] , GOUT[50] );
   BLOCK2 U351 (PIN[47] , PIN[49] , GIN[49] , GIN[51] , POUT[47] , GOUT[51] );
   BLOCK2 U352 (PIN[48] , PIN[50] , GIN[50] , GIN[52] , POUT[48] , GOUT[52] );
   BLOCK2 U353 (PIN[49] , PIN[51] , GIN[51] , GIN[53] , POUT[49] , GOUT[53] );
   BLOCK2 U354 (PIN[50] , PIN[52] , GIN[52] , GIN[54] , POUT[50] , GOUT[54] );
   BLOCK2 U355 (PIN[51] , PIN[53] , GIN[53] , GIN[55] , POUT[51] , GOUT[55] );
   BLOCK2 U356 (PIN[52] , PIN[54] , GIN[54] , GIN[56] , POUT[52] , GOUT[56] );
   BLOCK2 U357 (PIN[53] , PIN[55] , GIN[55] , GIN[57] , POUT[53] , GOUT[57] );
   BLOCK2 U358 (PIN[54] , PIN[56] , GIN[56] , GIN[58] , POUT[54] , GOUT[58] );
   BLOCK2 U359 (PIN[55] , PIN[57] , GIN[57] , GIN[59] , POUT[55] , GOUT[59] );
   BLOCK2 U360 (PIN[56] , PIN[58] , GIN[58] , GIN[60] , POUT[56] , GOUT[60] );
   BLOCK2 U361 (PIN[57] , PIN[59] , GIN[59] , GIN[61] , POUT[57] , GOUT[61] );
   BLOCK2 U362 (PIN[58] , PIN[60] , GIN[60] , GIN[62] , POUT[58] , GOUT[62] );
   BLOCK2 U363 (PIN[59] , PIN[61] , GIN[61] , GIN[63] , POUT[59] , GOUT[63] );
   BLOCK2 U364 (PIN[60] , PIN[62] , GIN[62] , GIN[64] , POUT[60] , GOUT[64] );
   
endmodule // DBLC_1_64


module DBLC_2_64 ( PIN, GIN, POUT, GOUT );
   
   input  [60:0] PIN;
   input [64:0]  GIN;
   
   output [56:0] POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   INVBLOCK U11 (GIN[1] , GOUT[1] );
   INVBLOCK U12 (GIN[2] , GOUT[2] );
   INVBLOCK U13 (GIN[3] , GOUT[3] );
   BLOCK1A U24 (PIN[0] , GIN[0] , GIN[4] , GOUT[4] );
   BLOCK1A U25 (PIN[1] , GIN[1] , GIN[5] , GOUT[5] );
   BLOCK1A U26 (PIN[2] , GIN[2] , GIN[6] , GOUT[6] );
   BLOCK1A U27 (PIN[3] , GIN[3] , GIN[7] , GOUT[7] );
   BLOCK1 U38 (PIN[0] , PIN[4] , GIN[4] , GIN[8] , POUT[0] , GOUT[8] );
   BLOCK1 U39 (PIN[1] , PIN[5] , GIN[5] , GIN[9] , POUT[1] , GOUT[9] );
   BLOCK1 U310 (PIN[2] , PIN[6] , GIN[6] , GIN[10] , POUT[2] , GOUT[10] );
   BLOCK1 U311 (PIN[3] , PIN[7] , GIN[7] , GIN[11] , POUT[3] , GOUT[11] );
   BLOCK1 U312 (PIN[4] , PIN[8] , GIN[8] , GIN[12] , POUT[4] , GOUT[12] );
   BLOCK1 U313 (PIN[5] , PIN[9] , GIN[9] , GIN[13] , POUT[5] , GOUT[13] );
   BLOCK1 U314 (PIN[6] , PIN[10] , GIN[10] , GIN[14] , POUT[6] , GOUT[14] );
   BLOCK1 U315 (PIN[7] , PIN[11] , GIN[11] , GIN[15] , POUT[7] , GOUT[15] );
   BLOCK1 U316 (PIN[8] , PIN[12] , GIN[12] , GIN[16] , POUT[8] , GOUT[16] );
   BLOCK1 U317 (PIN[9] , PIN[13] , GIN[13] , GIN[17] , POUT[9] , GOUT[17] );
   BLOCK1 U318 (PIN[10] , PIN[14] , GIN[14] , GIN[18] , POUT[10] , GOUT[18] );
   BLOCK1 U319 (PIN[11] , PIN[15] , GIN[15] , GIN[19] , POUT[11] , GOUT[19] );
   BLOCK1 U320 (PIN[12] , PIN[16] , GIN[16] , GIN[20] , POUT[12] , GOUT[20] );
   BLOCK1 U321 (PIN[13] , PIN[17] , GIN[17] , GIN[21] , POUT[13] , GOUT[21] );
   BLOCK1 U322 (PIN[14] , PIN[18] , GIN[18] , GIN[22] , POUT[14] , GOUT[22] );
   BLOCK1 U323 (PIN[15] , PIN[19] , GIN[19] , GIN[23] , POUT[15] , GOUT[23] );
   BLOCK1 U324 (PIN[16] , PIN[20] , GIN[20] , GIN[24] , POUT[16] , GOUT[24] );
   BLOCK1 U325 (PIN[17] , PIN[21] , GIN[21] , GIN[25] , POUT[17] , GOUT[25] );
   BLOCK1 U326 (PIN[18] , PIN[22] , GIN[22] , GIN[26] , POUT[18] , GOUT[26] );
   BLOCK1 U327 (PIN[19] , PIN[23] , GIN[23] , GIN[27] , POUT[19] , GOUT[27] );
   BLOCK1 U328 (PIN[20] , PIN[24] , GIN[24] , GIN[28] , POUT[20] , GOUT[28] );
   BLOCK1 U329 (PIN[21] , PIN[25] , GIN[25] , GIN[29] , POUT[21] , GOUT[29] );
   BLOCK1 U330 (PIN[22] , PIN[26] , GIN[26] , GIN[30] , POUT[22] , GOUT[30] );
   BLOCK1 U331 (PIN[23] , PIN[27] , GIN[27] , GIN[31] , POUT[23] , GOUT[31] );
   BLOCK1 U332 (PIN[24] , PIN[28] , GIN[28] , GIN[32] , POUT[24] , GOUT[32] );
   BLOCK1 U333 (PIN[25] , PIN[29] , GIN[29] , GIN[33] , POUT[25] , GOUT[33] );
   BLOCK1 U334 (PIN[26] , PIN[30] , GIN[30] , GIN[34] , POUT[26] , GOUT[34] );
   BLOCK1 U335 (PIN[27] , PIN[31] , GIN[31] , GIN[35] , POUT[27] , GOUT[35] );
   BLOCK1 U336 (PIN[28] , PIN[32] , GIN[32] , GIN[36] , POUT[28] , GOUT[36] );
   BLOCK1 U337 (PIN[29] , PIN[33] , GIN[33] , GIN[37] , POUT[29] , GOUT[37] );
   BLOCK1 U338 (PIN[30] , PIN[34] , GIN[34] , GIN[38] , POUT[30] , GOUT[38] );
   BLOCK1 U339 (PIN[31] , PIN[35] , GIN[35] , GIN[39] , POUT[31] , GOUT[39] );
   BLOCK1 U340 (PIN[32] , PIN[36] , GIN[36] , GIN[40] , POUT[32] , GOUT[40] );
   BLOCK1 U341 (PIN[33] , PIN[37] , GIN[37] , GIN[41] , POUT[33] , GOUT[41] );
   BLOCK1 U342 (PIN[34] , PIN[38] , GIN[38] , GIN[42] , POUT[34] , GOUT[42] );
   BLOCK1 U343 (PIN[35] , PIN[39] , GIN[39] , GIN[43] , POUT[35] , GOUT[43] );
   BLOCK1 U344 (PIN[36] , PIN[40] , GIN[40] , GIN[44] , POUT[36] , GOUT[44] );
   BLOCK1 U345 (PIN[37] , PIN[41] , GIN[41] , GIN[45] , POUT[37] , GOUT[45] );
   BLOCK1 U346 (PIN[38] , PIN[42] , GIN[42] , GIN[46] , POUT[38] , GOUT[46] );
   BLOCK1 U347 (PIN[39] , PIN[43] , GIN[43] , GIN[47] , POUT[39] , GOUT[47] );
   BLOCK1 U348 (PIN[40] , PIN[44] , GIN[44] , GIN[48] , POUT[40] , GOUT[48] );
   BLOCK1 U349 (PIN[41] , PIN[45] , GIN[45] , GIN[49] , POUT[41] , GOUT[49] );
   BLOCK1 U350 (PIN[42] , PIN[46] , GIN[46] , GIN[50] , POUT[42] , GOUT[50] );
   BLOCK1 U351 (PIN[43] , PIN[47] , GIN[47] , GIN[51] , POUT[43] , GOUT[51] );
   BLOCK1 U352 (PIN[44] , PIN[48] , GIN[48] , GIN[52] , POUT[44] , GOUT[52] );
   BLOCK1 U353 (PIN[45] , PIN[49] , GIN[49] , GIN[53] , POUT[45] , GOUT[53] );
   BLOCK1 U354 (PIN[46] , PIN[50] , GIN[50] , GIN[54] , POUT[46] , GOUT[54] );
   BLOCK1 U355 (PIN[47] , PIN[51] , GIN[51] , GIN[55] , POUT[47] , GOUT[55] );
   BLOCK1 U356 (PIN[48] , PIN[52] , GIN[52] , GIN[56] , POUT[48] , GOUT[56] );
   BLOCK1 U357 (PIN[49] , PIN[53] , GIN[53] , GIN[57] , POUT[49] , GOUT[57] );
   BLOCK1 U358 (PIN[50] , PIN[54] , GIN[54] , GIN[58] , POUT[50] , GOUT[58] );
   BLOCK1 U359 (PIN[51] , PIN[55] , GIN[55] , GIN[59] , POUT[51] , GOUT[59] );
   BLOCK1 U360 (PIN[52] , PIN[56] , GIN[56] , GIN[60] , POUT[52] , GOUT[60] );
   BLOCK1 U361 (PIN[53] , PIN[57] , GIN[57] , GIN[61] , POUT[53] , GOUT[61] );
   BLOCK1 U362 (PIN[54] , PIN[58] , GIN[58] , GIN[62] , POUT[54] , GOUT[62] );
   BLOCK1 U363 (PIN[55] , PIN[59] , GIN[59] , GIN[63] , POUT[55] , GOUT[63] );
   BLOCK1 U364 (PIN[56] , PIN[60] , GIN[60] , GIN[64] , POUT[56] , GOUT[64] );
   
endmodule // DBLC_2_64


module DBLC_3_64 ( PIN, GIN, POUT, GOUT );
   
   input  [56:0] PIN;
   input [64:0]  GIN;
   
   output [48:0] POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   INVBLOCK U11 (GIN[1] , GOUT[1] );
   INVBLOCK U12 (GIN[2] , GOUT[2] );
   INVBLOCK U13 (GIN[3] , GOUT[3] );
   INVBLOCK U14 (GIN[4] , GOUT[4] );
   INVBLOCK U15 (GIN[5] , GOUT[5] );
   INVBLOCK U16 (GIN[6] , GOUT[6] );
   INVBLOCK U17 (GIN[7] , GOUT[7] );
   BLOCK2A U28 (PIN[0] , GIN[0] , GIN[8] , GOUT[8] );
   BLOCK2A U29 (PIN[1] , GIN[1] , GIN[9] , GOUT[9] );
   BLOCK2A U210 (PIN[2] , GIN[2] , GIN[10] , GOUT[10] );
   BLOCK2A U211 (PIN[3] , GIN[3] , GIN[11] , GOUT[11] );
   BLOCK2A U212 (PIN[4] , GIN[4] , GIN[12] , GOUT[12] );
   BLOCK2A U213 (PIN[5] , GIN[5] , GIN[13] , GOUT[13] );
   BLOCK2A U214 (PIN[6] , GIN[6] , GIN[14] , GOUT[14] );
   BLOCK2A U215 (PIN[7] , GIN[7] , GIN[15] , GOUT[15] );
   BLOCK2 U316 (PIN[0] , PIN[8] , GIN[8] , GIN[16] , POUT[0] , GOUT[16] );
   BLOCK2 U317 (PIN[1] , PIN[9] , GIN[9] , GIN[17] , POUT[1] , GOUT[17] );
   BLOCK2 U318 (PIN[2] , PIN[10] , GIN[10] , GIN[18] , POUT[2] , GOUT[18] );
   BLOCK2 U319 (PIN[3] , PIN[11] , GIN[11] , GIN[19] , POUT[3] , GOUT[19] );
   BLOCK2 U320 (PIN[4] , PIN[12] , GIN[12] , GIN[20] , POUT[4] , GOUT[20] );
   BLOCK2 U321 (PIN[5] , PIN[13] , GIN[13] , GIN[21] , POUT[5] , GOUT[21] );
   BLOCK2 U322 (PIN[6] , PIN[14] , GIN[14] , GIN[22] , POUT[6] , GOUT[22] );
   BLOCK2 U323 (PIN[7] , PIN[15] , GIN[15] , GIN[23] , POUT[7] , GOUT[23] );
   BLOCK2 U324 (PIN[8] , PIN[16] , GIN[16] , GIN[24] , POUT[8] , GOUT[24] );
   BLOCK2 U325 (PIN[9] , PIN[17] , GIN[17] , GIN[25] , POUT[9] , GOUT[25] );
   BLOCK2 U326 (PIN[10] , PIN[18] , GIN[18] , GIN[26] , POUT[10] , GOUT[26] );
   BLOCK2 U327 (PIN[11] , PIN[19] , GIN[19] , GIN[27] , POUT[11] , GOUT[27] );
   BLOCK2 U328 (PIN[12] , PIN[20] , GIN[20] , GIN[28] , POUT[12] , GOUT[28] );
   BLOCK2 U329 (PIN[13] , PIN[21] , GIN[21] , GIN[29] , POUT[13] , GOUT[29] );
   BLOCK2 U330 (PIN[14] , PIN[22] , GIN[22] , GIN[30] , POUT[14] , GOUT[30] );
   BLOCK2 U331 (PIN[15] , PIN[23] , GIN[23] , GIN[31] , POUT[15] , GOUT[31] );
   BLOCK2 U332 (PIN[16] , PIN[24] , GIN[24] , GIN[32] , POUT[16] , GOUT[32] );
   BLOCK2 U333 (PIN[17] , PIN[25] , GIN[25] , GIN[33] , POUT[17] , GOUT[33] );
   BLOCK2 U334 (PIN[18] , PIN[26] , GIN[26] , GIN[34] , POUT[18] , GOUT[34] );
   BLOCK2 U335 (PIN[19] , PIN[27] , GIN[27] , GIN[35] , POUT[19] , GOUT[35] );
   BLOCK2 U336 (PIN[20] , PIN[28] , GIN[28] , GIN[36] , POUT[20] , GOUT[36] );
   BLOCK2 U337 (PIN[21] , PIN[29] , GIN[29] , GIN[37] , POUT[21] , GOUT[37] );
   BLOCK2 U338 (PIN[22] , PIN[30] , GIN[30] , GIN[38] , POUT[22] , GOUT[38] );
   BLOCK2 U339 (PIN[23] , PIN[31] , GIN[31] , GIN[39] , POUT[23] , GOUT[39] );
   BLOCK2 U340 (PIN[24] , PIN[32] , GIN[32] , GIN[40] , POUT[24] , GOUT[40] );
   BLOCK2 U341 (PIN[25] , PIN[33] , GIN[33] , GIN[41] , POUT[25] , GOUT[41] );
   BLOCK2 U342 (PIN[26] , PIN[34] , GIN[34] , GIN[42] , POUT[26] , GOUT[42] );
   BLOCK2 U343 (PIN[27] , PIN[35] , GIN[35] , GIN[43] , POUT[27] , GOUT[43] );
   BLOCK2 U344 (PIN[28] , PIN[36] , GIN[36] , GIN[44] , POUT[28] , GOUT[44] );
   BLOCK2 U345 (PIN[29] , PIN[37] , GIN[37] , GIN[45] , POUT[29] , GOUT[45] );
   BLOCK2 U346 (PIN[30] , PIN[38] , GIN[38] , GIN[46] , POUT[30] , GOUT[46] );
   BLOCK2 U347 (PIN[31] , PIN[39] , GIN[39] , GIN[47] , POUT[31] , GOUT[47] );
   BLOCK2 U348 (PIN[32] , PIN[40] , GIN[40] , GIN[48] , POUT[32] , GOUT[48] );
   BLOCK2 U349 (PIN[33] , PIN[41] , GIN[41] , GIN[49] , POUT[33] , GOUT[49] );
   BLOCK2 U350 (PIN[34] , PIN[42] , GIN[42] , GIN[50] , POUT[34] , GOUT[50] );
   BLOCK2 U351 (PIN[35] , PIN[43] , GIN[43] , GIN[51] , POUT[35] , GOUT[51] );
   BLOCK2 U352 (PIN[36] , PIN[44] , GIN[44] , GIN[52] , POUT[36] , GOUT[52] );
   BLOCK2 U353 (PIN[37] , PIN[45] , GIN[45] , GIN[53] , POUT[37] , GOUT[53] );
   BLOCK2 U354 (PIN[38] , PIN[46] , GIN[46] , GIN[54] , POUT[38] , GOUT[54] );
   BLOCK2 U355 (PIN[39] , PIN[47] , GIN[47] , GIN[55] , POUT[39] , GOUT[55] );
   BLOCK2 U356 (PIN[40] , PIN[48] , GIN[48] , GIN[56] , POUT[40] , GOUT[56] );
   BLOCK2 U357 (PIN[41] , PIN[49] , GIN[49] , GIN[57] , POUT[41] , GOUT[57] );
   BLOCK2 U358 (PIN[42] , PIN[50] , GIN[50] , GIN[58] , POUT[42] , GOUT[58] );
   BLOCK2 U359 (PIN[43] , PIN[51] , GIN[51] , GIN[59] , POUT[43] , GOUT[59] );
   BLOCK2 U360 (PIN[44] , PIN[52] , GIN[52] , GIN[60] , POUT[44] , GOUT[60] );
   BLOCK2 U361 (PIN[45] , PIN[53] , GIN[53] , GIN[61] , POUT[45] , GOUT[61] );
   BLOCK2 U362 (PIN[46] , PIN[54] , GIN[54] , GIN[62] , POUT[46] , GOUT[62] );
   BLOCK2 U363 (PIN[47] , PIN[55] , GIN[55] , GIN[63] , POUT[47] , GOUT[63] );
   BLOCK2 U364 (PIN[48] , PIN[56] , GIN[56] , GIN[64] , POUT[48] , GOUT[64] );
   
endmodule // DBLC_3_64


module DBLC_4_64 ( PIN, GIN, POUT, GOUT );
   
   input  [48:0] PIN;
   input [64:0]  GIN;
   
   output [32:0] POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   INVBLOCK U11 (GIN[1] , GOUT[1] );
   INVBLOCK U12 (GIN[2] , GOUT[2] );
   INVBLOCK U13 (GIN[3] , GOUT[3] );
   INVBLOCK U14 (GIN[4] , GOUT[4] );
   INVBLOCK U15 (GIN[5] , GOUT[5] );
   INVBLOCK U16 (GIN[6] , GOUT[6] );
   INVBLOCK U17 (GIN[7] , GOUT[7] );
   INVBLOCK U18 (GIN[8] , GOUT[8] );
   INVBLOCK U19 (GIN[9] , GOUT[9] );
   INVBLOCK U110 (GIN[10] , GOUT[10] );
   INVBLOCK U111 (GIN[11] , GOUT[11] );
   INVBLOCK U112 (GIN[12] , GOUT[12] );
   INVBLOCK U113 (GIN[13] , GOUT[13] );
   INVBLOCK U114 (GIN[14] , GOUT[14] );
   INVBLOCK U115 (GIN[15] , GOUT[15] );
   BLOCK1A U216 (PIN[0] , GIN[0] , GIN[16] , GOUT[16] );
   BLOCK1A U217 (PIN[1] , GIN[1] , GIN[17] , GOUT[17] );
   BLOCK1A U218 (PIN[2] , GIN[2] , GIN[18] , GOUT[18] );
   BLOCK1A U219 (PIN[3] , GIN[3] , GIN[19] , GOUT[19] );
   BLOCK1A U220 (PIN[4] , GIN[4] , GIN[20] , GOUT[20] );
   BLOCK1A U221 (PIN[5] , GIN[5] , GIN[21] , GOUT[21] );
   BLOCK1A U222 (PIN[6] , GIN[6] , GIN[22] , GOUT[22] );
   BLOCK1A U223 (PIN[7] , GIN[7] , GIN[23] , GOUT[23] );
   BLOCK1A U224 (PIN[8] , GIN[8] , GIN[24] , GOUT[24] );
   BLOCK1A U225 (PIN[9] , GIN[9] , GIN[25] , GOUT[25] );
   BLOCK1A U226 (PIN[10] , GIN[10] , GIN[26] , GOUT[26] );
   BLOCK1A U227 (PIN[11] , GIN[11] , GIN[27] , GOUT[27] );
   BLOCK1A U228 (PIN[12] , GIN[12] , GIN[28] , GOUT[28] );
   BLOCK1A U229 (PIN[13] , GIN[13] , GIN[29] , GOUT[29] );
   BLOCK1A U230 (PIN[14] , GIN[14] , GIN[30] , GOUT[30] );
   BLOCK1A U231 (PIN[15] , GIN[15] , GIN[31] , GOUT[31] );
   BLOCK1 U332 (PIN[0] , PIN[16] , GIN[16] , GIN[32] , POUT[0] , GOUT[32] );
   BLOCK1 U333 (PIN[1] , PIN[17] , GIN[17] , GIN[33] , POUT[1] , GOUT[33] );
   BLOCK1 U334 (PIN[2] , PIN[18] , GIN[18] , GIN[34] , POUT[2] , GOUT[34] );
   BLOCK1 U335 (PIN[3] , PIN[19] , GIN[19] , GIN[35] , POUT[3] , GOUT[35] );
   BLOCK1 U336 (PIN[4] , PIN[20] , GIN[20] , GIN[36] , POUT[4] , GOUT[36] );
   BLOCK1 U337 (PIN[5] , PIN[21] , GIN[21] , GIN[37] , POUT[5] , GOUT[37] );
   BLOCK1 U338 (PIN[6] , PIN[22] , GIN[22] , GIN[38] , POUT[6] , GOUT[38] );
   BLOCK1 U339 (PIN[7] , PIN[23] , GIN[23] , GIN[39] , POUT[7] , GOUT[39] );
   BLOCK1 U340 (PIN[8] , PIN[24] , GIN[24] , GIN[40] , POUT[8] , GOUT[40] );
   BLOCK1 U341 (PIN[9] , PIN[25] , GIN[25] , GIN[41] , POUT[9] , GOUT[41] );
   BLOCK1 U342 (PIN[10] , PIN[26] , GIN[26] , GIN[42] , POUT[10] , GOUT[42] );
   BLOCK1 U343 (PIN[11] , PIN[27] , GIN[27] , GIN[43] , POUT[11] , GOUT[43] );
   BLOCK1 U344 (PIN[12] , PIN[28] , GIN[28] , GIN[44] , POUT[12] , GOUT[44] );
   BLOCK1 U345 (PIN[13] , PIN[29] , GIN[29] , GIN[45] , POUT[13] , GOUT[45] );
   BLOCK1 U346 (PIN[14] , PIN[30] , GIN[30] , GIN[46] , POUT[14] , GOUT[46] );
   BLOCK1 U347 (PIN[15] , PIN[31] , GIN[31] , GIN[47] , POUT[15] , GOUT[47] );
   BLOCK1 U348 (PIN[16] , PIN[32] , GIN[32] , GIN[48] , POUT[16] , GOUT[48] );
   BLOCK1 U349 (PIN[17] , PIN[33] , GIN[33] , GIN[49] , POUT[17] , GOUT[49] );
   BLOCK1 U350 (PIN[18] , PIN[34] , GIN[34] , GIN[50] , POUT[18] , GOUT[50] );
   BLOCK1 U351 (PIN[19] , PIN[35] , GIN[35] , GIN[51] , POUT[19] , GOUT[51] );
   BLOCK1 U352 (PIN[20] , PIN[36] , GIN[36] , GIN[52] , POUT[20] , GOUT[52] );
   BLOCK1 U353 (PIN[21] , PIN[37] , GIN[37] , GIN[53] , POUT[21] , GOUT[53] );
   BLOCK1 U354 (PIN[22] , PIN[38] , GIN[38] , GIN[54] , POUT[22] , GOUT[54] );
   BLOCK1 U355 (PIN[23] , PIN[39] , GIN[39] , GIN[55] , POUT[23] , GOUT[55] );
   BLOCK1 U356 (PIN[24] , PIN[40] , GIN[40] , GIN[56] , POUT[24] , GOUT[56] );
   BLOCK1 U357 (PIN[25] , PIN[41] , GIN[41] , GIN[57] , POUT[25] , GOUT[57] );
   BLOCK1 U358 (PIN[26] , PIN[42] , GIN[42] , GIN[58] , POUT[26] , GOUT[58] );
   BLOCK1 U359 (PIN[27] , PIN[43] , GIN[43] , GIN[59] , POUT[27] , GOUT[59] );
   BLOCK1 U360 (PIN[28] , PIN[44] , GIN[44] , GIN[60] , POUT[28] , GOUT[60] );
   BLOCK1 U361 (PIN[29] , PIN[45] , GIN[45] , GIN[61] , POUT[29] , GOUT[61] );
   BLOCK1 U362 (PIN[30] , PIN[46] , GIN[46] , GIN[62] , POUT[30] , GOUT[62] );
   BLOCK1 U363 (PIN[31] , PIN[47] , GIN[47] , GIN[63] , POUT[31] , GOUT[63] );
   BLOCK1 U364 (PIN[32] , PIN[48] , GIN[48] , GIN[64] , POUT[32] , GOUT[64] );
   
endmodule // DBLC_4_64


module DBLC_5_64 ( PIN, GIN, POUT, GOUT );
   
   input  [32:0] PIN;
   input [64:0]  GIN;
   
   output [0:0]  POUT;
   output [64:0] GOUT;
   
   INVBLOCK U10 (GIN[0] , GOUT[0] );
   INVBLOCK U11 (GIN[1] , GOUT[1] );
   INVBLOCK U12 (GIN[2] , GOUT[2] );
   INVBLOCK U13 (GIN[3] , GOUT[3] );
   INVBLOCK U14 (GIN[4] , GOUT[4] );
   INVBLOCK U15 (GIN[5] , GOUT[5] );
   INVBLOCK U16 (GIN[6] , GOUT[6] );
   INVBLOCK U17 (GIN[7] , GOUT[7] );
   INVBLOCK U18 (GIN[8] , GOUT[8] );
   INVBLOCK U19 (GIN[9] , GOUT[9] );
   INVBLOCK U110 (GIN[10] , GOUT[10] );
   INVBLOCK U111 (GIN[11] , GOUT[11] );
   INVBLOCK U112 (GIN[12] , GOUT[12] );
   INVBLOCK U113 (GIN[13] , GOUT[13] );
   INVBLOCK U114 (GIN[14] , GOUT[14] );
   INVBLOCK U115 (GIN[15] , GOUT[15] );
   INVBLOCK U116 (GIN[16] , GOUT[16] );
   INVBLOCK U117 (GIN[17] , GOUT[17] );
   INVBLOCK U118 (GIN[18] , GOUT[18] );
   INVBLOCK U119 (GIN[19] , GOUT[19] );
   INVBLOCK U120 (GIN[20] , GOUT[20] );
   INVBLOCK U121 (GIN[21] , GOUT[21] );
   INVBLOCK U122 (GIN[22] , GOUT[22] );
   INVBLOCK U123 (GIN[23] , GOUT[23] );
   INVBLOCK U124 (GIN[24] , GOUT[24] );
   INVBLOCK U125 (GIN[25] , GOUT[25] );
   INVBLOCK U126 (GIN[26] , GOUT[26] );
   INVBLOCK U127 (GIN[27] , GOUT[27] );
   INVBLOCK U128 (GIN[28] , GOUT[28] );
   INVBLOCK U129 (GIN[29] , GOUT[29] );
   INVBLOCK U130 (GIN[30] , GOUT[30] );
   INVBLOCK U131 (GIN[31] , GOUT[31] );
   BLOCK2A U232 (PIN[0] , GIN[0] , GIN[32] , GOUT[32] );
   BLOCK2A U233 (PIN[1] , GIN[1] , GIN[33] , GOUT[33] );
   BLOCK2A U234 (PIN[2] , GIN[2] , GIN[34] , GOUT[34] );
   BLOCK2A U235 (PIN[3] , GIN[3] , GIN[35] , GOUT[35] );
   BLOCK2A U236 (PIN[4] , GIN[4] , GIN[36] , GOUT[36] );
   BLOCK2A U237 (PIN[5] , GIN[5] , GIN[37] , GOUT[37] );
   BLOCK2A U238 (PIN[6] , GIN[6] , GIN[38] , GOUT[38] );
   BLOCK2A U239 (PIN[7] , GIN[7] , GIN[39] , GOUT[39] );
   BLOCK2A U240 (PIN[8] , GIN[8] , GIN[40] , GOUT[40] );
   BLOCK2A U241 (PIN[9] , GIN[9] , GIN[41] , GOUT[41] );
   BLOCK2A U242 (PIN[10] , GIN[10] , GIN[42] , GOUT[42] );
   BLOCK2A U243 (PIN[11] , GIN[11] , GIN[43] , GOUT[43] );
   BLOCK2A U244 (PIN[12] , GIN[12] , GIN[44] , GOUT[44] );
   BLOCK2A U245 (PIN[13] , GIN[13] , GIN[45] , GOUT[45] );
   BLOCK2A U246 (PIN[14] , GIN[14] , GIN[46] , GOUT[46] );
   BLOCK2A U247 (PIN[15] , GIN[15] , GIN[47] , GOUT[47] );
   BLOCK2A U248 (PIN[16] , GIN[16] , GIN[48] , GOUT[48] );
   BLOCK2A U249 (PIN[17] , GIN[17] , GIN[49] , GOUT[49] );
   BLOCK2A U250 (PIN[18] , GIN[18] , GIN[50] , GOUT[50] );
   BLOCK2A U251 (PIN[19] , GIN[19] , GIN[51] , GOUT[51] );
   BLOCK2A U252 (PIN[20] , GIN[20] , GIN[52] , GOUT[52] );
   BLOCK2A U253 (PIN[21] , GIN[21] , GIN[53] , GOUT[53] );
   BLOCK2A U254 (PIN[22] , GIN[22] , GIN[54] , GOUT[54] );
   BLOCK2A U255 (PIN[23] , GIN[23] , GIN[55] , GOUT[55] );
   BLOCK2A U256 (PIN[24] , GIN[24] , GIN[56] , GOUT[56] );
   BLOCK2A U257 (PIN[25] , GIN[25] , GIN[57] , GOUT[57] );
   BLOCK2A U258 (PIN[26] , GIN[26] , GIN[58] , GOUT[58] );
   BLOCK2A U259 (PIN[27] , GIN[27] , GIN[59] , GOUT[59] );
   BLOCK2A U260 (PIN[28] , GIN[28] , GIN[60] , GOUT[60] );
   BLOCK2A U261 (PIN[29] , GIN[29] , GIN[61] , GOUT[61] );
   BLOCK2A U262 (PIN[30] , GIN[30] , GIN[62] , GOUT[62] );
   BLOCK2A U263 (PIN[31] , GIN[31] , GIN[63] , GOUT[63] );
   BLOCK2 U364 (PIN[0] , PIN[32] , GIN[32] , GIN[64] , POUT[0] , GOUT[64] );
   
endmodule // DBLC_5_64


module XORSTAGE_64 ( A, B, PBIT, CARRY, SUM, COUT );
   
   input  [63:0] A;
   input [63:0]  B;
   input 	 PBIT;
   input [64:0]  CARRY;
   
   output [63:0] SUM;
   output 	 COUT;
   
   XXOR1 U20 (A[0] , B[0] , CARRY[0] , SUM[0] );
   XXOR1 U21 (A[1] , B[1] , CARRY[1] , SUM[1] );
   XXOR1 U22 (A[2] , B[2] , CARRY[2] , SUM[2] );
   XXOR1 U23 (A[3] , B[3] , CARRY[3] , SUM[3] );
   XXOR1 U24 (A[4] , B[4] , CARRY[4] , SUM[4] );
   XXOR1 U25 (A[5] , B[5] , CARRY[5] , SUM[5] );
   XXOR1 U26 (A[6] , B[6] , CARRY[6] , SUM[6] );
   XXOR1 U27 (A[7] , B[7] , CARRY[7] , SUM[7] );
   XXOR1 U28 (A[8] , B[8] , CARRY[8] , SUM[8] );
   XXOR1 U29 (A[9] , B[9] , CARRY[9] , SUM[9] );
   XXOR1 U210 (A[10] , B[10] , CARRY[10] , SUM[10] );
   XXOR1 U211 (A[11] , B[11] , CARRY[11] , SUM[11] );
   XXOR1 U212 (A[12] , B[12] , CARRY[12] , SUM[12] );
   XXOR1 U213 (A[13] , B[13] , CARRY[13] , SUM[13] );
   XXOR1 U214 (A[14] , B[14] , CARRY[14] , SUM[14] );
   XXOR1 U215 (A[15] , B[15] , CARRY[15] , SUM[15] );
   XXOR1 U216 (A[16] , B[16] , CARRY[16] , SUM[16] );
   XXOR1 U217 (A[17] , B[17] , CARRY[17] , SUM[17] );
   XXOR1 U218 (A[18] , B[18] , CARRY[18] , SUM[18] );
   XXOR1 U219 (A[19] , B[19] , CARRY[19] , SUM[19] );
   XXOR1 U220 (A[20] , B[20] , CARRY[20] , SUM[20] );
   XXOR1 U221 (A[21] , B[21] , CARRY[21] , SUM[21] );
   XXOR1 U222 (A[22] , B[22] , CARRY[22] , SUM[22] );
   XXOR1 U223 (A[23] , B[23] , CARRY[23] , SUM[23] );
   XXOR1 U224 (A[24] , B[24] , CARRY[24] , SUM[24] );
   XXOR1 U225 (A[25] , B[25] , CARRY[25] , SUM[25] );
   XXOR1 U226 (A[26] , B[26] , CARRY[26] , SUM[26] );
   XXOR1 U227 (A[27] , B[27] , CARRY[27] , SUM[27] );
   XXOR1 U228 (A[28] , B[28] , CARRY[28] , SUM[28] );
   XXOR1 U229 (A[29] , B[29] , CARRY[29] , SUM[29] );
   XXOR1 U230 (A[30] , B[30] , CARRY[30] , SUM[30] );
   XXOR1 U231 (A[31] , B[31] , CARRY[31] , SUM[31] );
   XXOR1 U232 (A[32] , B[32] , CARRY[32] , SUM[32] );
   XXOR1 U233 (A[33] , B[33] , CARRY[33] , SUM[33] );
   XXOR1 U234 (A[34] , B[34] , CARRY[34] , SUM[34] );
   XXOR1 U235 (A[35] , B[35] , CARRY[35] , SUM[35] );
   XXOR1 U236 (A[36] , B[36] , CARRY[36] , SUM[36] );
   XXOR1 U237 (A[37] , B[37] , CARRY[37] , SUM[37] );
   XXOR1 U238 (A[38] , B[38] , CARRY[38] , SUM[38] );
   XXOR1 U239 (A[39] , B[39] , CARRY[39] , SUM[39] );
   XXOR1 U240 (A[40] , B[40] , CARRY[40] , SUM[40] );
   XXOR1 U241 (A[41] , B[41] , CARRY[41] , SUM[41] );
   XXOR1 U242 (A[42] , B[42] , CARRY[42] , SUM[42] );
   XXOR1 U243 (A[43] , B[43] , CARRY[43] , SUM[43] );
   XXOR1 U244 (A[44] , B[44] , CARRY[44] , SUM[44] );
   XXOR1 U245 (A[45] , B[45] , CARRY[45] , SUM[45] );
   XXOR1 U246 (A[46] , B[46] , CARRY[46] , SUM[46] );
   XXOR1 U247 (A[47] , B[47] , CARRY[47] , SUM[47] );
   XXOR1 U248 (A[48] , B[48] , CARRY[48] , SUM[48] );
   XXOR1 U249 (A[49] , B[49] , CARRY[49] , SUM[49] );
   XXOR1 U250 (A[50] , B[50] , CARRY[50] , SUM[50] );
   XXOR1 U251 (A[51] , B[51] , CARRY[51] , SUM[51] );
   XXOR1 U252 (A[52] , B[52] , CARRY[52] , SUM[52] );
   XXOR1 U253 (A[53] , B[53] , CARRY[53] , SUM[53] );
   XXOR1 U254 (A[54] , B[54] , CARRY[54] , SUM[54] );
   XXOR1 U255 (A[55] , B[55] , CARRY[55] , SUM[55] );
   XXOR1 U256 (A[56] , B[56] , CARRY[56] , SUM[56] );
   XXOR1 U257 (A[57] , B[57] , CARRY[57] , SUM[57] );
   XXOR1 U258 (A[58] , B[58] , CARRY[58] , SUM[58] );
   XXOR1 U259 (A[59] , B[59] , CARRY[59] , SUM[59] );
   XXOR1 U260 (A[60] , B[60] , CARRY[60] , SUM[60] );
   XXOR1 U261 (A[61] , B[61] , CARRY[61] , SUM[61] );
   XXOR1 U262 (A[62] , B[62] , CARRY[62] , SUM[62] );
   XXOR1 U263 (A[63] , B[63] , CARRY[63] , SUM[63] );
   BLOCK1A U1 (PBIT , CARRY[0] , CARRY[64] , COUT );
   
endmodule // XORSTAGE_64


module DBLCTREE_64 ( PIN, GIN, GOUT, POUT );
   
   input  [63:0] PIN;
   input [64:0]  GIN;
   
   output [64:0] GOUT;
   output [0:0]  POUT;
   
   wire [62:0] 	 INTPROP_0;
   wire [64:0] 	 INTGEN_0;
   wire [60:0] 	 INTPROP_1;
   wire [64:0] 	 INTGEN_1;
   wire [56:0] 	 INTPROP_2;
   wire [64:0] 	 INTGEN_2;
   wire [48:0] 	 INTPROP_3;
   wire [64:0] 	 INTGEN_3;
   wire [32:0] 	 INTPROP_4;
   wire [64:0] 	 INTGEN_4;
   
   DBLC_0_64 U_0 (.PIN(PIN) , .GIN(GIN) , .POUT(INTPROP_0) , .GOUT(INTGEN_0) );
   DBLC_1_64 U_1 (.PIN(INTPROP_0) , .GIN(INTGEN_0) , .POUT(INTPROP_1) , .GOUT(INTGEN_1) );
   DBLC_2_64 U_2 (.PIN(INTPROP_1) , .GIN(INTGEN_1) , .POUT(INTPROP_2) , .GOUT(INTGEN_2) );
   DBLC_3_64 U_3 (.PIN(INTPROP_2) , .GIN(INTGEN_2) , .POUT(INTPROP_3) , .GOUT(INTGEN_3) );
   DBLC_4_64 U_4 (.PIN(INTPROP_3) , .GIN(INTGEN_3) , .POUT(INTPROP_4) , .GOUT(INTGEN_4) );
   DBLC_5_64 U_5 (.PIN(INTPROP_4) , .GIN(INTGEN_4) , .POUT(POUT) , .GOUT(GOUT) );
   
endmodule // DBLCTREE_64


module DBLCADDER_64_64 ( OPA, OPB, CIN, SUM, COUT );
   
   input  [63:0] OPA;
   input [63:0]  OPB;
   input 	 CIN;
   
   output [63:0] SUM;
   output 	 COUT;
   
   wire [63:0] 	 INTPROP;
   wire [64:0] 	 INTGEN;
   wire [0:0] 	 PBIT;
   wire [64:0] 	 CARRY;
   
   PRESTAGE_64 U1 (OPA , OPB , CIN , INTPROP , INTGEN );
   DBLCTREE_64 U2 (INTPROP , INTGEN , CARRY , PBIT );
   XORSTAGE_64 U3 (OPA[63:0] , OPB[63:0] , PBIT[0] , CARRY[64:0] , SUM , COUT );
   
endmodule 

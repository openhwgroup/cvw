///////////////////////////////////////////
//
// Written: me@KatherineParry.com
// Modified: 7/5/2022
//
// Purpose: Leading Zero Counter
// 
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////
//leading zero counter i.e. priority encoder
module lzc #(parameter WIDTH = 1) (
    input logic  [WIDTH-1:0]            num,
    output logic [$clog2(WIDTH+1)-1:0]  ZeroCnt
);
/* verilator lint_off CMPCONST */
/* verilator lint_off WIDTH */
    
    logic [31:0] i;
    always_comb begin
        i = 0;
        while (~num[WIDTH-1-i] & (i < WIDTH)) i = i+1;  // search for leading one
        ZeroCnt = i;
    end
/* verilator lint_on WIDTH */
/* verilator lint_on CMPCONST */
endmodule

localparam VPN_SEGMENT_BITS = (LLEN == 32 ? 10 : 9);


 parameter cvw_t P = '{ 
    PA_BITS : PA_BITS,
    XLEN:     XLEN,
    AHBW:     AHBW,
    MISA:     MISA,
    BUS_SUPPORTED: BUS_SUPPORTED,
    ZICSR_SUPPORTED: ZICSR_SUPPORTED,
    M_SUPPORTED: M_SUPPORTED,
    ZMMUL_SUPPORTED: ZMMUL_SUPPORTED,
    F_SUPPORTED: F_SUPPORTED,
    PMP_ENTRIES: PMP_ENTRIES,
    LLEN:     LLEN,
    FPGA:     FPGA,
    QEMU:     QEMU,
    VPN_SEGMENT_BITS: VPN_SEGMENT_BITS,
   FLEN:     FLEN
};
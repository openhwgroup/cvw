///////////////////////////////////////////
// tests.vh
//
// Written: David_Harris@hmc.edu 7 October 2021
// Modified: 
//
// Purpose: List of tests to apply
// 
// A component of the Wally configurable RISC-V project.
// 
// Copyright (C) 2021 Harvey Mudd College & Oklahoma State University
//
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, 
// modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software 
// is furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES 
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS 
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT 
// OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
///////////////////////////////////////////

`define IMPERASTEST   "0"
`define RISCVARCHTEST "1"
`define WALLYTEST "2"
`define MYIMPERASTEST   "3"
`define COREMARK "4"
`define EMBENCH "5"
// *** remove MYIMPERASTEST cases when ported 

string tvpaths[] = '{
    "../../addins/imperas-riscv-tests/work/",
    "../../tests/riscof/work/",
    "../../tests/wally-riscv-arch-test/work/",
    "../../tests/imperas-riscv-tests/work/",
    "../../benchmarks/riscv-coremark/work/",
    "../../addins/embench-iot/bd_speed/src/"
};

  string coremark[] = '{
    `COREMARK,
    "coremark.bare.riscv"
  };

  string embench[] = '{
    `EMBENCH,
    "aha-mont64/aha-mont64",
    "crc32/crc32",
    "cubic/cubic",
    "edn/edn",
    "huffbench/huffbench",
    "matmult-int/matmult-int",
    "md5sum/md5sum",
    "minver/minver",
    "nbody/nbody",
    "nettle-aes/nettle-aes",
    "nettle-sha256/nettle-sha256",
    "nsichneu/nsichneu",
    "picojpeg/picojpeg",
    "primecount/primecount",
    "qrduino/qrduino",
    "sglib-combined/sglib-combined",
    "slre/slre",
    "st/st",
    "statemate/statemate",
    "tarfind/tarfind",
    "ud/ud",
    "wikisort/wikisort"
  };

  string wally64a[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-amo",
    "rv64i_m/privilege/WALLY-lrsc",
    "rv64i_m/privilege/WALLY-status-fp-enabled-01"
  };

    string wally32a[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/WALLY-amo",
    "rv32i_m/privilege/WALLY-lrsc",
    "rv32i_m/privilege/WALLY-status-fp-enabled-01"

  };

  // *** restore CSR tests from Imperas old

    string extra64i[] = '{
    `MYIMPERASTEST,
    "rv64i_m/I/WALLY-ADD",
    "rv64i_m/I/WALLY-SUB",
    "rv64i_m/I/WALLY-ADDI",
    "rv64i_m/I/WALLY-ANDI",
    "rv64i_m/I/WALLY-ORI",
    "rv64i_m/I/WALLY-XORI",
    "rv64i_m/I/WALLY-SLTI",
    "rv64i_m/I/WALLY-SLTIU",
    "rv64i_m/I/WALLY-SLLI",
    "rv64i_m/I/WALLY-SRLI",
    "rv64i_m/I/WALLY-SRAI",
    "rv64i_m/I/WALLY-JAL",
    "rv64i_m/I/WALLY-JALR",
    "rv64i_m/I/WALLY-STORE",
    "rv64i_m/I/WALLY-ADDIW",
    "rv64i_m/I/WALLY-SLLIW",
    "rv64i_m/I/WALLY-SRLIW",
    "rv64i_m/I/WALLY-SRAIW",
    "rv64i_m/I/WALLY-ADDW",
    "rv64i_m/I/WALLY-SUBW",
    "rv64i_m/I/WALLY-SLLW",
    "rv64i_m/I/WALLY-SRLW",
    "rv64i_m/I/WALLY-SRAW",
    "rv64i_m/I/WALLY-BEQ",
    "rv64i_m/I/WALLY-BNE",
    "rv64i_m/I/WALLY-BLTU",
    "rv64i_m/I/WALLY-BLT",
    "rv64i_m/I/WALLY-BGE",
    "rv64i_m/I/WALLY-BGEU",
    "rv64i_m/I/WALLY-CSRRW",
    "rv64i_m/I/WALLY-CSRRS",
    "rv64i_m/I/WALLY-CSRRC",
    "rv64i_m/I/WALLY-CSRRWI",
    "rv64i_m/I/WALLY-CSRRSI",
    "rv64i_m/I/WALLY-CSRRCI" 
  };

  
string imperas32f[] = '{
    `IMPERASTEST,
    "rv32i_m/F/FADD-S-DYN-RDN-01",
    "rv32i_m/F/FADD-S-DYN-RMM-01",
    "rv32i_m/F/FADD-S-DYN-RNE-01",
    "rv32i_m/F/FADD-S-DYN-RTZ-01",
    "rv32i_m/F/FADD-S-DYN-RUP-01",
    "rv32i_m/F/FADD-S-RDN-01",
    "rv32i_m/F/FADD-S-RMM-01",
    "rv32i_m/F/FADD-S-RNE-01",
    "rv32i_m/F/FADD-S-RTZ-01",
    "rv32i_m/F/FADD-S-RUP-01",
    "rv32i_m/F/FCLASS-S-01",
    "rv32i_m/F/FCVT-S-W-DYN-RDN-01",
    "rv32i_m/F/FCVT-S-W-DYN-RMM-01",
    "rv32i_m/F/FCVT-S-W-DYN-RNE-01",
    "rv32i_m/F/FCVT-S-W-DYN-RTZ-01",
    "rv32i_m/F/FCVT-S-W-DYN-RUP-01",
    "rv32i_m/F/FCVT-S-W-RDN-01",
    "rv32i_m/F/FCVT-S-W-RMM-01",
    "rv32i_m/F/FCVT-S-W-RNE-01",
    "rv32i_m/F/FCVT-S-W-RTZ-01",
    "rv32i_m/F/FCVT-S-W-RUP-01",
    "rv32i_m/F/FCVT-S-WU-DYN-RDN-01",
    "rv32i_m/F/FCVT-S-WU-DYN-RMM-01",
    "rv32i_m/F/FCVT-S-WU-DYN-RNE-01",
    "rv32i_m/F/FCVT-S-WU-DYN-RTZ-01",
    "rv32i_m/F/FCVT-S-WU-DYN-RUP-01",
    "rv32i_m/F/FCVT-S-WU-RDN-01",
    "rv32i_m/F/FCVT-S-WU-RMM-01",
    "rv32i_m/F/FCVT-S-WU-RNE-01",
    "rv32i_m/F/FCVT-S-WU-RTZ-01",
    "rv32i_m/F/FCVT-S-WU-RUP-01",
    "rv32i_m/F/FCVT-W-S-DYN-RDN-01",
    "rv32i_m/F/FCVT-W-S-DYN-RMM-01",
    "rv32i_m/F/FCVT-W-S-DYN-RNE-01",
    "rv32i_m/F/FCVT-W-S-DYN-RTZ-01",
    "rv32i_m/F/FCVT-W-S-DYN-RUP-01",
    "rv32i_m/F/FCVT-W-S-RDN-01",
    "rv32i_m/F/FCVT-W-S-RMM-01",
    "rv32i_m/F/FCVT-W-S-RNE-01",
    "rv32i_m/F/FCVT-W-S-RTZ-01",
    "rv32i_m/F/FCVT-W-S-RUP-01",
    "rv32i_m/F/FCVT-WU-S-DYN-RDN-01",
    "rv32i_m/F/FCVT-WU-S-DYN-RMM-01",
    "rv32i_m/F/FCVT-WU-S-DYN-RNE-01",
    "rv32i_m/F/FCVT-WU-S-DYN-RTZ-01",
    "rv32i_m/F/FCVT-WU-S-DYN-RUP-01",
    "rv32i_m/F/FCVT-WU-S-RDN-01",
    "rv32i_m/F/FCVT-WU-S-RMM-01",
    "rv32i_m/F/FCVT-WU-S-RNE-01",
    "rv32i_m/F/FCVT-WU-S-RTZ-01",
    "rv32i_m/F/FCVT-WU-S-RUP-01",
    // "rv32i_m/F/FDIV-S-DYN-RDN-01",
    // "rv32i_m/F/FDIV-S-DYN-RMM-01",
    // "rv32i_m/F/FDIV-S-DYN-RNE-01",
    // "rv32i_m/F/FDIV-S-DYN-RTZ-01",
    // "rv32i_m/F/FDIV-S-DYN-RUP-01",
    // "rv32i_m/F/FDIV-S-RDN-01",
    // "rv32i_m/F/FDIV-S-RMM-01",
    // "rv32i_m/F/FDIV-S-RNE-01",
    // "rv32i_m/F/FDIV-S-RTZ-01",
    // "rv32i_m/F/FDIV-S-RUP-01",
    "rv32i_m/F/FEQ-S-01",
    "rv32i_m/F/FLE-S-01",
    "rv32i_m/F/FLT-S-01",
    "rv32i_m/F/FLW-01",
    "rv32i_m/F/FMADD-S-DYN-RDN-01",
    "rv32i_m/F/FMADD-S-DYN-RMM-01",
    "rv32i_m/F/FMADD-S-DYN-RNE-01",
    "rv32i_m/F/FMADD-S-DYN-RTZ-01",
    "rv32i_m/F/FMADD-S-DYN-RUP-01",
    "rv32i_m/F/FMADD-S-RDN-01",
    "rv32i_m/F/FMADD-S-RMM-01",
    "rv32i_m/F/FMADD-S-RNE-01",
    "rv32i_m/F/FMADD-S-RTZ-01",
    "rv32i_m/F/FMADD-S-RUP-01",
    "rv32i_m/F/FMAX-S-01",
    "rv32i_m/F/FMIN-S-01",
    "rv32i_m/F/FMSUB-S-DYN-RDN-01",
    "rv32i_m/F/FMSUB-S-DYN-RMM-01",
    "rv32i_m/F/FMSUB-S-DYN-RNE-01",
    "rv32i_m/F/FMSUB-S-DYN-RTZ-01",
    "rv32i_m/F/FMSUB-S-DYN-RUP-01",
    "rv32i_m/F/FMSUB-S-RDN-01",
    "rv32i_m/F/FMSUB-S-RMM-01",
    "rv32i_m/F/FMSUB-S-RNE-01",
    "rv32i_m/F/FMSUB-S-RTZ-01",
    "rv32i_m/F/FMSUB-S-RUP-01",
    "rv32i_m/F/FMUL-S-DYN-RDN-01",
    "rv32i_m/F/FMUL-S-DYN-RMM-01",
    "rv32i_m/F/FMUL-S-DYN-RNE-01",
    "rv32i_m/F/FMUL-S-DYN-RTZ-01",
    "rv32i_m/F/FMUL-S-DYN-RUP-01",
    "rv32i_m/F/FMUL-S-RDN-01",
    "rv32i_m/F/FMUL-S-RMM-01",
    "rv32i_m/F/FMUL-S-RNE-01",
    "rv32i_m/F/FMUL-S-RTZ-01",
    "rv32i_m/F/FMUL-S-RUP-01",
    "rv32i_m/F/FMV-W-X-01",
    "rv32i_m/F/FMV-X-W-01",
    "rv32i_m/F/FNMADD-S-DYN-RDN-01",
    "rv32i_m/F/FNMADD-S-DYN-RMM-01",
    "rv32i_m/F/FNMADD-S-DYN-RNE-01",
    "rv32i_m/F/FNMADD-S-DYN-RTZ-01",
    "rv32i_m/F/FNMADD-S-DYN-RUP-01",
    "rv32i_m/F/FNMADD-S-RDN-01",
    "rv32i_m/F/FNMADD-S-RMM-01",
    "rv32i_m/F/FNMADD-S-RNE-01",
    "rv32i_m/F/FNMADD-S-RTZ-01",
    "rv32i_m/F/FNMADD-S-RUP-01",
    "rv32i_m/F/FNMSUB-S-DYN-RDN-01",
    "rv32i_m/F/FNMSUB-S-DYN-RMM-01",
    "rv32i_m/F/FNMSUB-S-DYN-RNE-01",
    "rv32i_m/F/FNMSUB-S-DYN-RTZ-01",
    "rv32i_m/F/FNMSUB-S-DYN-RUP-01",
    "rv32i_m/F/FNMSUB-S-RDN-01",
    "rv32i_m/F/FNMSUB-S-RMM-01",
    "rv32i_m/F/FNMSUB-S-RNE-01",
    "rv32i_m/F/FNMSUB-S-RTZ-01",
    "rv32i_m/F/FNMSUB-S-RUP-01",
    "rv32i_m/F/FSGNJN-S-01",
    "rv32i_m/F/FSGNJ-S-01",
    "rv32i_m/F/FSGNJX-S-01",
    // "rv32i_m/F/FSQRT-S-DYN-RDN-01",
    // "rv32i_m/F/FSQRT-S-DYN-RMM-01",
    // "rv32i_m/F/FSQRT-S-DYN-RNE-01",
    // "rv32i_m/F/FSQRT-S-DYN-RTZ-01",
    // "rv32i_m/F/FSQRT-S-DYN-RUP-01",
    // "rv32i_m/F/FSQRT-S-RDN-01",
    // "rv32i_m/F/FSQRT-S-RMM-01",
    // "rv32i_m/F/FSQRT-S-RNE-01",
    // "rv32i_m/F/FSQRT-S-RTZ-01",
    // "rv32i_m/F/FSQRT-S-RUP-01",
    "rv32i_m/F/FSUB-S-DYN-RDN-01",
    "rv32i_m/F/FSUB-S-DYN-RMM-01",
    "rv32i_m/F/FSUB-S-DYN-RNE-01",
    "rv32i_m/F/FSUB-S-DYN-RTZ-01",
    "rv32i_m/F/FSUB-S-DYN-RUP-01",
    "rv32i_m/F/FSUB-S-RDN-01",
    "rv32i_m/F/FSUB-S-RMM-01",
    "rv32i_m/F/FSUB-S-RNE-01",
    "rv32i_m/F/FSUB-S-RTZ-01",
    "rv32i_m/F/FSUB-S-RUP-01",
    "rv32i_m/F/FSW-01"
  };

  string imperas64f[] = '{
    `IMPERASTEST,
    "rv64i_m/F/FADD-S-DYN-RDN-01",
    "rv64i_m/F/FADD-S-DYN-RMM-01",
    "rv64i_m/F/FADD-S-DYN-RNE-01",
    "rv64i_m/F/FADD-S-DYN-RTZ-01",
    "rv64i_m/F/FADD-S-DYN-RUP-01",
    "rv64i_m/F/FADD-S-RDN-01",
    "rv64i_m/F/FADD-S-RMM-01",
    "rv64i_m/F/FADD-S-RNE-01",
    "rv64i_m/F/FADD-S-RTZ-01",
    "rv64i_m/F/FADD-S-RUP-01",
    "rv64i_m/F/FCLASS-S-01",
    "rv64i_m/F/FCVT-L-S-DYN-RDN-01",
    "rv64i_m/F/FCVT-L-S-DYN-RMM-01",
    "rv64i_m/F/FCVT-L-S-DYN-RNE-01",
    "rv64i_m/F/FCVT-L-S-DYN-RTZ-01",
    "rv64i_m/F/FCVT-L-S-DYN-RUP-01",
    "rv64i_m/F/FCVT-L-S-RDN-01",
    "rv64i_m/F/FCVT-L-S-RMM-01",
    "rv64i_m/F/FCVT-L-S-RNE-01",
    "rv64i_m/F/FCVT-L-S-RTZ-01",
    "rv64i_m/F/FCVT-L-S-RUP-01",
    "rv64i_m/F/FCVT-LU-S-DYN-RDN-01",
    "rv64i_m/F/FCVT-LU-S-DYN-RMM-01",
    "rv64i_m/F/FCVT-LU-S-DYN-RNE-01",
    "rv64i_m/F/FCVT-LU-S-DYN-RTZ-01",
    "rv64i_m/F/FCVT-LU-S-DYN-RUP-01",
    "rv64i_m/F/FCVT-LU-S-RDN-01",
    "rv64i_m/F/FCVT-LU-S-RMM-01",
    "rv64i_m/F/FCVT-LU-S-RNE-01",
    "rv64i_m/F/FCVT-LU-S-RTZ-01",
    "rv64i_m/F/FCVT-LU-S-RUP-01",
    "rv64i_m/F/FCVT-S-L-DYN-RDN-01",
    "rv64i_m/F/FCVT-S-L-DYN-RMM-01",
    "rv64i_m/F/FCVT-S-L-DYN-RNE-01",
    "rv64i_m/F/FCVT-S-L-DYN-RTZ-01",
    "rv64i_m/F/FCVT-S-L-DYN-RUP-01",
    "rv64i_m/F/FCVT-S-L-RDN-01",
    "rv64i_m/F/FCVT-S-L-RMM-01",
    "rv64i_m/F/FCVT-S-L-RNE-01",
    "rv64i_m/F/FCVT-S-L-RTZ-01",
    "rv64i_m/F/FCVT-S-L-RUP-01",
    "rv64i_m/F/FCVT-S-LU-DYN-RDN-01",
    "rv64i_m/F/FCVT-S-LU-DYN-RMM-01",
    "rv64i_m/F/FCVT-S-LU-DYN-RNE-01",
    "rv64i_m/F/FCVT-S-LU-DYN-RTZ-01",
    "rv64i_m/F/FCVT-S-LU-DYN-RUP-01",
    "rv64i_m/F/FCVT-S-LU-RDN-01",
    "rv64i_m/F/FCVT-S-LU-RMM-01",
    "rv64i_m/F/FCVT-S-LU-RNE-01",
    "rv64i_m/F/FCVT-S-LU-RTZ-01",
    "rv64i_m/F/FCVT-S-LU-RUP-01",
    "rv64i_m/F/FCVT-S-W-DYN-RDN-01",
    "rv64i_m/F/FCVT-S-W-DYN-RMM-01",
    "rv64i_m/F/FCVT-S-W-DYN-RNE-01",
    "rv64i_m/F/FCVT-S-W-DYN-RTZ-01",
    "rv64i_m/F/FCVT-S-W-DYN-RUP-01",
    "rv64i_m/F/FCVT-S-W-RDN-01",
    "rv64i_m/F/FCVT-S-W-RMM-01",
    "rv64i_m/F/FCVT-S-W-RNE-01",
    "rv64i_m/F/FCVT-S-W-RTZ-01",
    "rv64i_m/F/FCVT-S-W-RUP-01",
    "rv64i_m/F/FCVT-S-WU-DYN-RDN-01",
    "rv64i_m/F/FCVT-S-WU-DYN-RMM-01",
    "rv64i_m/F/FCVT-S-WU-DYN-RNE-01",
    "rv64i_m/F/FCVT-S-WU-DYN-RTZ-01",
    "rv64i_m/F/FCVT-S-WU-DYN-RUP-01",
    "rv64i_m/F/FCVT-S-WU-RDN-01",
    "rv64i_m/F/FCVT-S-WU-RMM-01",
    "rv64i_m/F/FCVT-S-WU-RNE-01",
    "rv64i_m/F/FCVT-S-WU-RTZ-01",
    "rv64i_m/F/FCVT-S-WU-RUP-01",
    "rv64i_m/F/FCVT-W-S-DYN-RDN-01",
    "rv64i_m/F/FCVT-W-S-DYN-RMM-01",
    "rv64i_m/F/FCVT-W-S-DYN-RNE-01",
    "rv64i_m/F/FCVT-W-S-DYN-RTZ-01",
    "rv64i_m/F/FCVT-W-S-DYN-RUP-01",
    "rv64i_m/F/FCVT-W-S-RDN-01",
    "rv64i_m/F/FCVT-W-S-RMM-01",
    "rv64i_m/F/FCVT-W-S-RNE-01",
    "rv64i_m/F/FCVT-W-S-RTZ-01",
    "rv64i_m/F/FCVT-W-S-RUP-01",
    "rv64i_m/F/FCVT-WU-S-DYN-RDN-01",
    "rv64i_m/F/FCVT-WU-S-DYN-RMM-01",
    "rv64i_m/F/FCVT-WU-S-DYN-RNE-01",
    "rv64i_m/F/FCVT-WU-S-DYN-RTZ-01",
    "rv64i_m/F/FCVT-WU-S-DYN-RUP-01",
    "rv64i_m/F/FCVT-WU-S-RDN-01",
    "rv64i_m/F/FCVT-WU-S-RMM-01",
    "rv64i_m/F/FCVT-WU-S-RNE-01",
    "rv64i_m/F/FCVT-WU-S-RTZ-01",
    "rv64i_m/F/FCVT-WU-S-RUP-01",
    // "rv64i_m/F/FDIV-S-DYN-RDN-01",
    // "rv64i_m/F/FDIV-S-DYN-RMM-01",
    // "rv64i_m/F/FDIV-S-DYN-RNE-01",
    // "rv64i_m/F/FDIV-S-DYN-RTZ-01",
    // "rv64i_m/F/FDIV-S-DYN-RUP-01",
    // "rv64i_m/F/FDIV-S-RDN-01",
    // "rv64i_m/F/FDIV-S-RMM-01",
    // "rv64i_m/F/FDIV-S-RNE-01",
    // "rv64i_m/F/FDIV-S-RTZ-01",
    // "rv64i_m/F/FDIV-S-RUP-01",
    "rv64i_m/F/FEQ-S-01",
    "rv64i_m/F/FLE-S-01",
    "rv64i_m/F/FLT-S-01",
    "rv64i_m/F/FLW-01",
    "rv64i_m/F/FMADD-S-DYN-RDN-01",
    "rv64i_m/F/FMADD-S-DYN-RMM-01",
    "rv64i_m/F/FMADD-S-DYN-RNE-01",
    "rv64i_m/F/FMADD-S-DYN-RTZ-01",
    "rv64i_m/F/FMADD-S-DYN-RUP-01",
    "rv64i_m/F/FMADD-S-RDN-01",
    "rv64i_m/F/FMADD-S-RMM-01",
    "rv64i_m/F/FMADD-S-RNE-01",
    "rv64i_m/F/FMADD-S-RTZ-01",
    "rv64i_m/F/FMADD-S-RUP-01",
    "rv64i_m/F/FMAX-S-01",
    "rv64i_m/F/FMIN-S-01",
    "rv64i_m/F/FMSUB-S-DYN-RDN-01",
    "rv64i_m/F/FMSUB-S-DYN-RMM-01",
    "rv64i_m/F/FMSUB-S-DYN-RNE-01",
    "rv64i_m/F/FMSUB-S-DYN-RTZ-01",
    "rv64i_m/F/FMSUB-S-DYN-RUP-01",
    "rv64i_m/F/FMSUB-S-RDN-01",
    "rv64i_m/F/FMSUB-S-RMM-01",
    "rv64i_m/F/FMSUB-S-RNE-01",
    "rv64i_m/F/FMSUB-S-RTZ-01",
    "rv64i_m/F/FMSUB-S-RUP-01",
    "rv64i_m/F/FMUL-S-DYN-RDN-01",
    "rv64i_m/F/FMUL-S-DYN-RMM-01",
    "rv64i_m/F/FMUL-S-DYN-RNE-01",
    "rv64i_m/F/FMUL-S-DYN-RTZ-01",
    "rv64i_m/F/FMUL-S-DYN-RUP-01",
    "rv64i_m/F/FMUL-S-RDN-01",
    "rv64i_m/F/FMUL-S-RMM-01",
    "rv64i_m/F/FMUL-S-RNE-01",
    "rv64i_m/F/FMUL-S-RTZ-01",
    "rv64i_m/F/FMUL-S-RUP-01",
    "rv64i_m/F/FMV-W-X-01",
    "rv64i_m/F/FMV-X-W-01",
    "rv64i_m/F/FNMADD-S-DYN-RDN-01",
    "rv64i_m/F/FNMADD-S-DYN-RMM-01",
    "rv64i_m/F/FNMADD-S-DYN-RNE-01",
    "rv64i_m/F/FNMADD-S-DYN-RTZ-01",
    "rv64i_m/F/FNMADD-S-DYN-RUP-01",
    "rv64i_m/F/FNMADD-S-RDN-01",
    "rv64i_m/F/FNMADD-S-RMM-01",
    "rv64i_m/F/FNMADD-S-RNE-01",
    "rv64i_m/F/FNMADD-S-RTZ-01",
    "rv64i_m/F/FNMADD-S-RUP-01",
    "rv64i_m/F/FNMSUB-S-DYN-RDN-01",
    "rv64i_m/F/FNMSUB-S-DYN-RMM-01",
    "rv64i_m/F/FNMSUB-S-DYN-RNE-01",
    "rv64i_m/F/FNMSUB-S-DYN-RTZ-01",
    "rv64i_m/F/FNMSUB-S-DYN-RUP-01",
    "rv64i_m/F/FNMSUB-S-RDN-01",
    "rv64i_m/F/FNMSUB-S-RMM-01",
    "rv64i_m/F/FNMSUB-S-RNE-01",
    "rv64i_m/F/FNMSUB-S-RTZ-01",
    "rv64i_m/F/FNMSUB-S-RUP-01",
    "rv64i_m/F/FSGNJN-S-01",
    "rv64i_m/F/FSGNJ-S-01",
    "rv64i_m/F/FSGNJX-S-01",
    // "rv64i_m/F/FSQRT-S-DYN-RDN-01",
    // "rv64i_m/F/FSQRT-S-DYN-RMM-01",
    // "rv64i_m/F/FSQRT-S-DYN-RNE-01",
    // "rv64i_m/F/FSQRT-S-DYN-RTZ-01",
    // "rv64i_m/F/FSQRT-S-DYN-RUP-01",
    // "rv64i_m/F/FSQRT-S-RDN-01",
    // "rv64i_m/F/FSQRT-S-RMM-01",
    // "rv64i_m/F/FSQRT-S-RNE-01",
    // "rv64i_m/F/FSQRT-S-RTZ-01",
    // "rv64i_m/F/FSQRT-S-RUP-01",
    "rv64i_m/F/FSUB-S-DYN-RDN-01",
    "rv64i_m/F/FSUB-S-DYN-RMM-01",
    "rv64i_m/F/FSUB-S-DYN-RNE-01",
    "rv64i_m/F/FSUB-S-DYN-RTZ-01",
    "rv64i_m/F/FSUB-S-DYN-RUP-01",
    "rv64i_m/F/FSUB-S-RDN-01",
    "rv64i_m/F/FSUB-S-RMM-01",
    "rv64i_m/F/FSUB-S-RNE-01",
    "rv64i_m/F/FSUB-S-RTZ-01",
    "rv64i_m/F/FSUB-S-RUP-01",
    "rv64i_m/F/FSW-01"
  };

  string imperas64d[] = '{
    `IMPERASTEST,
    "rv64i_m/D/FADD-D-DYN-RDN-01",
    "rv64i_m/D/FADD-D-DYN-RMM-01",
    "rv64i_m/D/FADD-D-DYN-RNE-01",
    "rv64i_m/D/FADD-D-DYN-RTZ-01",
    "rv64i_m/D/FADD-D-DYN-RUP-01",
    "rv64i_m/D/FADD-D-RDN-01",
    "rv64i_m/D/FADD-D-RMM-01",
    "rv64i_m/D/FADD-D-RNE-01",
    "rv64i_m/D/FADD-D-RTZ-01",
    "rv64i_m/D/FADD-D-RUP-01",
    "rv64i_m/D/FCLASS-D-01",
    "rv64i_m/D/FCVT-D-L-DYN-RDN-01",
    "rv64i_m/D/FCVT-D-L-DYN-RMM-01",
    "rv64i_m/D/FCVT-D-L-DYN-RNE-01",
    "rv64i_m/D/FCVT-D-L-DYN-RTZ-01",
    "rv64i_m/D/FCVT-D-L-DYN-RUP-01",
    "rv64i_m/D/FCVT-D-L-RDN-01",
    "rv64i_m/D/FCVT-D-L-RMM-01",
    "rv64i_m/D/FCVT-D-L-RNE-01",
    "rv64i_m/D/FCVT-D-L-RTZ-01",
    "rv64i_m/D/FCVT-D-L-RUP-01",
    "rv64i_m/D/FCVT-D-LU-DYN-RDN-01",
    "rv64i_m/D/FCVT-D-LU-DYN-RMM-01",
    "rv64i_m/D/FCVT-D-LU-DYN-RNE-01",
    "rv64i_m/D/FCVT-D-LU-DYN-RTZ-01",
    "rv64i_m/D/FCVT-D-LU-DYN-RUP-01",
    "rv64i_m/D/FCVT-D-LU-RDN-01",
    "rv64i_m/D/FCVT-D-LU-RMM-01",
    "rv64i_m/D/FCVT-D-LU-RNE-01",
    "rv64i_m/D/FCVT-D-LU-RTZ-01",
    "rv64i_m/D/FCVT-D-LU-RUP-01",
    "rv64i_m/D/FCVT-D-S-01",
    "rv64i_m/D/FCVT-D-W-01",
    "rv64i_m/D/FCVT-D-WU-01",
    "rv64i_m/D/FCVT-L-D-DYN-RDN-01",
    "rv64i_m/D/FCVT-L-D-DYN-RMM-01",
    "rv64i_m/D/FCVT-L-D-DYN-RNE-01",
    "rv64i_m/D/FCVT-L-D-DYN-RTZ-01",
    "rv64i_m/D/FCVT-L-D-DYN-RUP-01",
    "rv64i_m/D/FCVT-L-D-RDN-01",
    "rv64i_m/D/FCVT-L-D-RMM-01",
    "rv64i_m/D/FCVT-L-D-RNE-01",
    "rv64i_m/D/FCVT-L-D-RTZ-01",
    "rv64i_m/D/FCVT-L-D-RUP-01",
    "rv64i_m/D/FCVT-LU-D-DYN-RDN-01",
    "rv64i_m/D/FCVT-LU-D-DYN-RMM-01",
    "rv64i_m/D/FCVT-LU-D-DYN-RNE-01",
    "rv64i_m/D/FCVT-LU-D-DYN-RTZ-01",
    "rv64i_m/D/FCVT-LU-D-DYN-RUP-01",
    "rv64i_m/D/FCVT-LU-D-RDN-01",
    "rv64i_m/D/FCVT-LU-D-RMM-01",
    "rv64i_m/D/FCVT-LU-D-RNE-01",
    "rv64i_m/D/FCVT-LU-D-RTZ-01",
    "rv64i_m/D/FCVT-LU-D-RUP-01",
    "rv64i_m/D/FCVT-S-D-DYN-RDN-01",
    "rv64i_m/D/FCVT-S-D-DYN-RMM-01",
    "rv64i_m/D/FCVT-S-D-DYN-RNE-01",
    "rv64i_m/D/FCVT-S-D-DYN-RTZ-01",
    "rv64i_m/D/FCVT-S-D-DYN-RUP-01",
    "rv64i_m/D/FCVT-S-D-RDN-01",
    "rv64i_m/D/FCVT-S-D-RMM-01",
    "rv64i_m/D/FCVT-S-D-RNE-01",
    "rv64i_m/D/FCVT-S-D-RTZ-01",
    "rv64i_m/D/FCVT-S-D-RUP-01",
    "rv64i_m/D/FCVT-W-D-DYN-RDN-01",
    "rv64i_m/D/FCVT-W-D-DYN-RMM-01",
    "rv64i_m/D/FCVT-W-D-DYN-RNE-01",
    "rv64i_m/D/FCVT-W-D-DYN-RTZ-01",
    "rv64i_m/D/FCVT-W-D-DYN-RUP-01",
    "rv64i_m/D/FCVT-W-D-RDN-01",
    "rv64i_m/D/FCVT-W-D-RMM-01",
    "rv64i_m/D/FCVT-W-D-RNE-01",
    "rv64i_m/D/FCVT-W-D-RTZ-01",
    "rv64i_m/D/FCVT-W-D-RUP-01",
    "rv64i_m/D/FCVT-WU-D-DYN-RDN-01",
    "rv64i_m/D/FCVT-WU-D-DYN-RMM-01",
    "rv64i_m/D/FCVT-WU-D-DYN-RNE-01",
    "rv64i_m/D/FCVT-WU-D-DYN-RTZ-01",
    "rv64i_m/D/FCVT-WU-D-DYN-RUP-01",
    "rv64i_m/D/FCVT-WU-D-RDN-01",
    "rv64i_m/D/FCVT-WU-D-RMM-01",
    "rv64i_m/D/FCVT-WU-D-RNE-01",
    "rv64i_m/D/FCVT-WU-D-RTZ-01",
    "rv64i_m/D/FCVT-WU-D-RUP-01",
    // "rv64i_m/D/FDIV-D-DYN-RDN-01",
    // "rv64i_m/D/FDIV-D-DYN-RMM-01",
    // "rv64i_m/D/FDIV-D-DYN-RNE-01",
    // "rv64i_m/D/FDIV-D-DYN-RTZ-01",
    // "rv64i_m/D/FDIV-D-DYN-RUP-01",
    // "rv64i_m/D/FDIV-D-RDN-01",
    // "rv64i_m/D/FDIV-D-RMM-01",
    // "rv64i_m/D/FDIV-D-RNE-01",
    // "rv64i_m/D/FDIV-D-RTZ-01",
    // "rv64i_m/D/FDIV-D-RUP-01",
    "rv64i_m/D/FEQ-D-01",
    "rv64i_m/D/FLD-01",
    "rv64i_m/D/FLE-D-01",
    "rv64i_m/D/FLT-D-01",
    "rv64i_m/D/FMADD-D-DYN-RDN-01",
    "rv64i_m/D/FMADD-D-DYN-RMM-01",
    "rv64i_m/D/FMADD-D-DYN-RNE-01",
    "rv64i_m/D/FMADD-D-DYN-RTZ-01",
    "rv64i_m/D/FMADD-D-DYN-RUP-01",
    "rv64i_m/D/FMADD-D-RDN-01",
    "rv64i_m/D/FMADD-D-RMM-01",
    "rv64i_m/D/FMADD-D-RNE-01",
    "rv64i_m/D/FMADD-D-RTZ-01",
    "rv64i_m/D/FMADD-D-RUP-01",
    "rv64i_m/D/FMAX-D-01",
    "rv64i_m/D/FMIN-D-01",
    "rv64i_m/D/FMSUB-D-DYN-RDN-01",
    "rv64i_m/D/FMSUB-D-DYN-RMM-01",
    "rv64i_m/D/FMSUB-D-DYN-RNE-01",
    "rv64i_m/D/FMSUB-D-DYN-RTZ-01",
    "rv64i_m/D/FMSUB-D-DYN-RUP-01",
    "rv64i_m/D/FMSUB-D-RDN-01",
    "rv64i_m/D/FMSUB-D-RMM-01",
    "rv64i_m/D/FMSUB-D-RNE-01",
    "rv64i_m/D/FMSUB-D-RTZ-01",
    "rv64i_m/D/FMSUB-D-RUP-01",
    "rv64i_m/D/FMUL-D-DYN-RDN-01",
    "rv64i_m/D/FMUL-D-DYN-RMM-01",
    "rv64i_m/D/FMUL-D-DYN-RNE-01",
    "rv64i_m/D/FMUL-D-DYN-RTZ-01",
    "rv64i_m/D/FMUL-D-DYN-RUP-01",
    "rv64i_m/D/FMUL-D-RDN-01",
    "rv64i_m/D/FMUL-D-RMM-01",
    "rv64i_m/D/FMUL-D-RNE-01",
    "rv64i_m/D/FMUL-D-RTZ-01",
    "rv64i_m/D/FMUL-D-RUP-01",
    "rv64i_m/D/FMV-D-X-01",
    "rv64i_m/D/FMV-X-D-01",
    "rv64i_m/D/FNMADD-D-DYN-RDN-01",
    "rv64i_m/D/FNMADD-D-DYN-RMM-01",
    "rv64i_m/D/FNMADD-D-DYN-RNE-01",
    "rv64i_m/D/FNMADD-D-DYN-RTZ-01",
    "rv64i_m/D/FNMADD-D-DYN-RUP-01",
    "rv64i_m/D/FNMADD-D-RDN-01",
    "rv64i_m/D/FNMADD-D-RMM-01",
    "rv64i_m/D/FNMADD-D-RNE-01",
    "rv64i_m/D/FNMADD-D-RTZ-01",
    "rv64i_m/D/FNMADD-D-RUP-01",
    "rv64i_m/D/FNMSUB-D-DYN-RDN-01",
    "rv64i_m/D/FNMSUB-D-DYN-RMM-01",
    "rv64i_m/D/FNMSUB-D-DYN-RNE-01",
    "rv64i_m/D/FNMSUB-D-DYN-RTZ-01",
    "rv64i_m/D/FNMSUB-D-DYN-RUP-01",
    "rv64i_m/D/FNMSUB-D-RDN-01",
    "rv64i_m/D/FNMSUB-D-RMM-01",
    "rv64i_m/D/FNMSUB-D-RNE-01",
    "rv64i_m/D/FNMSUB-D-RTZ-01",
    "rv64i_m/D/FNMSUB-D-RUP-01",
    "rv64i_m/D/FSD-01",
    "rv64i_m/D/FSGNJ-D-01",
    "rv64i_m/D/FSGNJN-D-01",
    "rv64i_m/D/FSGNJX-D-01",
    // "rv64i_m/D/FSQRT-D-DYN-RDN-01",
    // "rv64i_m/D/FSQRT-D-DYN-RMM-01",
    // "rv64i_m/D/FSQRT-D-DYN-RNE-01",
    // "rv64i_m/D/FSQRT-D-DYN-RTZ-01",
    // "rv64i_m/D/FSQRT-D-DYN-RUP-01",
    // "rv64i_m/D/FSQRT-D-RDN-01",
    // "rv64i_m/D/FSQRT-D-RMM-01",
    // "rv64i_m/D/FSQRT-D-RNE-01",
    // "rv64i_m/D/FSQRT-D-RTZ-01",
    // "rv64i_m/D/FSQRT-D-RUP-01",
    "rv64i_m/D/FSUB-D-DYN-RDN-01",
    "rv64i_m/D/FSUB-D-DYN-RMM-01",
    "rv64i_m/D/FSUB-D-DYN-RNE-01",
    "rv64i_m/D/FSUB-D-DYN-RTZ-01",
    "rv64i_m/D/FSUB-D-DYN-RUP-01",
    "rv64i_m/D/FSUB-D-RDN-01",
    "rv64i_m/D/FSUB-D-RMM-01",
    "rv64i_m/D/FSUB-D-RNE-01",
    "rv64i_m/D/FSUB-D-RTZ-01",
    "rv64i_m/D/FSUB-D-RUP-01"
};

  string imperas64m[] = '{
    `IMPERASTEST,
    "rv64i_m/M/DIV-01",
    "rv64i_m/M/DIVU-01",
    "rv64i_m/M/DIVUW-01",
    "rv64i_m/M/DIVW-01",
    "rv64i_m/M/MUL-01",
    "rv64i_m/M/MULH-01",
    "rv64i_m/M/MULHSU-01",
    "rv64i_m/M/MULHU-01",
    "rv64i_m/M/MULW-01",
    "rv64i_m/M/REM-01",
    "rv64i_m/M/REMU-01",
    "rv64i_m/M/REMUW-01",
    "rv64i_m/M/REMW-01"
  };

  string imperas64c[] = '{
    `IMPERASTEST,
    "rv64i_m/C/C-ADD-01",
    "rv64i_m/C/C-ADDI-01",
    "rv64i_m/C/C-ADDI16SP-01",
    "rv64i_m/C/C-ADDI4SPN-01",
    "rv64i_m/C/C-ADDIW-01",
    "rv64i_m/C/C-ADDW-01",
    "rv64i_m/C/C-AND-01",
    "rv64i_m/C/C-ANDI-01",
    "rv64i_m/C/C-BEQZ-01",
    "rv64i_m/C/C-BNEZ-01",
    "rv64i_m/C/C-J-01",
    "rv64i_m/C/C-JALR-01",
    "rv64i_m/C/C-JR-01",
    "rv64i_m/C/C-LD-01",
    "rv64i_m/C/C-LDSP-01",
    "rv64i_m/C/C-LI-01",
    "rv64i_m/C/C-LUI-01",
    "rv64i_m/C/C-LW-01",
    "rv64i_m/C/C-LWSP-01",
    "rv64i_m/C/C-MV-01",
    "rv64i_m/C/C-OR-01",
    "rv64i_m/C/C-SD-01",
    "rv64i_m/C/C-SDSP-01",
    "rv64i_m/C/C-SLLI-01",
    "rv64i_m/C/C-SRAI-01",
    "rv64i_m/C/C-SRLI-01",
    "rv64i_m/C/C-SUB-01",
    "rv64i_m/C/C-SUBW-01",
    "rv64i_m/C/C-SW-01",
    "rv64i_m/C/C-SWSP-01",
    "rv64i_m/C/C-XOR-01",
    "rv64i_m/C/I-C-EBREAK-01",
    "rv64i_m/C/I-C-NOP-01"
  };

  string imperas64iNOc[] = {
    `IMPERASTEST,
    "rv64i_m/I/I-MISALIGN_JMP-01"
  };

  string imperas64i[] = '{
    `IMPERASTEST,
    "rv64i_m/I/I-DELAY_SLOTS-01",
    "rv64i_m/I/ADD-01",
    "rv64i_m/I/ADDI-01",
    "rv64i_m/I/ADDIW-01",
    "rv64i_m/I/ADDW-01",
    "rv64i_m/I/AND-01",
    "rv64i_m/I/ANDI-01",
    "rv64i_m/I/AUIPC-01",
    "rv64i_m/I/BEQ-01",
    "rv64i_m/I/BGE-01",
    "rv64i_m/I/BGEU-01",
    "rv64i_m/I/BLT-01",
    "rv64i_m/I/BLTU-01",
    "rv64i_m/I/BNE-01",
    "rv64i_m/I/I-DELAY_SLOTS-01",
    "rv64i_m/I/I-EBREAK-01",
    "rv64i_m/I/I-ECALL-01",
    "rv64i_m/I/I-ENDIANESS-01",
    "rv64i_m/I/I-IO-01",
//    "rv64i_m/I/I-MISALIGN_JMP-01",
    "rv64i_m/I/I-MISALIGN_LDST-01",
    "rv64i_m/I/I-NOP-01",
    "rv64i_m/I/I-RF_size-01",
    "rv64i_m/I/I-RF_width-01",
    "rv64i_m/I/I-RF_x0-01",
    "rv64i_m/I/JAL-01",
    "rv64i_m/I/JALR-01",
    "rv64i_m/I/LB-01",
    "rv64i_m/I/LBU-01",
    "rv64i_m/I/LD-01",
    "rv64i_m/I/LH-01",
    "rv64i_m/I/LHU-01",
    "rv64i_m/I/LUI-01",
    "rv64i_m/I/LW-01",
    "rv64i_m/I/LWU-01",
    "rv64i_m/I/OR-01",
    "rv64i_m/I/ORI-01",
    "rv64i_m/I/SB-01",
    "rv64i_m/I/SD-01",
    "rv64i_m/I/SH-01",
    "rv64i_m/I/SLL-01",
    "rv64i_m/I/SLLI-01",
    "rv64i_m/I/SLLIW-01",
    "rv64i_m/I/SLLW-01",
    "rv64i_m/I/SLT-01",
    "rv64i_m/I/SLTI-01",
    "rv64i_m/I/SLTIU-01",
    "rv64i_m/I/SLTU-01",
    "rv64i_m/I/SRA-01",
    "rv64i_m/I/SRAI-01",
    "rv64i_m/I/SRAIW-01",
    "rv64i_m/I/SRAW-01",
    "rv64i_m/I/SRL-01",
    "rv64i_m/I/SRLI-01",
    "rv64i_m/I/SRLIW-01",
    "rv64i_m/I/SRLW-01",
    "rv64i_m/I/SUB-01",
    "rv64i_m/I/SUBW-01",
    "rv64i_m/I/SW-01",
    "rv64i_m/I/XOR-01",
    "rv64i_m/I/XORI-01"
  };

  string imperas32m[] = '{
    `IMPERASTEST,
    "rv32i_m/M/DIV-01",
    "rv32i_m/M/DIVU-01",
    "rv32i_m/M/MUL-01",
    "rv32i_m/M/MULH-01",
    "rv32i_m/M/MULHSU-01",
    "rv32i_m/M/MULHU-01",
    "rv32i_m/M/REM-01",
    "rv32i_m/M/REMU-01"
  };

  string imperas32c[] = '{
    `IMPERASTEST,
    "rv32i_m/C/C-ADD-01",
    "rv32i_m/C/C-ADDI-01",
    "rv32i_m/C/C-ADDI16SP-01",
    "rv32i_m/C/C-ADDI4SPN-01",
    "rv32i_m/C/C-AND-01",
    "rv32i_m/C/C-ANDI-01",
    "rv32i_m/C/C-BEQZ-01",
    "rv32i_m/C/C-BNEZ-01",
    "rv32i_m/C/C-J-01",
    "rv32i_m/C/C-JAL-01",
    "rv32i_m/C/C-JALR-01",
    "rv32i_m/C/C-JR-01",
    "rv32i_m/C/C-LI-01",
    "rv32i_m/C/C-LUI-01",
    "rv32i_m/C/C-LW-01",
    "rv32i_m/C/C-LWSP-01",
    "rv32i_m/C/C-MV-01",
    "rv32i_m/C/C-OR-01",
    "rv32i_m/C/C-SLLI-01",
    "rv32i_m/C/C-SRAI-01",
    "rv32i_m/C/C-SRLI-01",
    "rv32i_m/C/C-SUB-01",
    "rv32i_m/C/C-SW-01",
    "rv32i_m/C/C-SWSP-01",
    "rv32i_m/C/C-XOR-01",
    "rv32i_m/C/I-C-EBREAK-01",
    "rv32i_m/C/I-C-NOP-01"
  };

  string imperas32iNOc[] = {
    `IMPERASTEST,
    "rv32i_m/I/I-MISALIGN_JMP-01"
  };

  string imperas32i[] = {
    `IMPERASTEST,
    "rv32i_m/I/ADD-01",
    "rv32i_m/I/ADDI-01",
    "rv32i_m/I/AND-01",
    "rv32i_m/I/ANDI-01",
    "rv32i_m/I/AUIPC-01",
    "rv32i_m/I/BEQ-01",
    "rv32i_m/I/BGE-01",
    "rv32i_m/I/BGEU-01",
    "rv32i_m/I/BLT-01",
    "rv32i_m/I/BLTU-01",
    "rv32i_m/I/BNE-01",
    "rv32i_m/I/I-DELAY_SLOTS-01",
    "rv32i_m/I/I-EBREAK-01",
    "rv32i_m/I/I-ECALL-01",
    "rv32i_m/I/I-ENDIANESS-01",
    "rv32i_m/I/I-IO-01",
//    "rv32i_m/I/I-MISALIGN_JMP-01",
    "rv32i_m/I/I-MISALIGN_LDST-01",
    "rv32i_m/I/I-NOP-01",
    "rv32i_m/I/I-RF_size-01",
    "rv32i_m/I/I-RF_width-01",
    "rv32i_m/I/I-RF_x0-01",
    "rv32i_m/I/JAL-01",
    "rv32i_m/I/JALR-01",
    "rv32i_m/I/LB-01",
    "rv32i_m/I/LBU-01",
    "rv32i_m/I/LH-01",
    "rv32i_m/I/LHU-01",
    "rv32i_m/I/LUI-01",
    "rv32i_m/I/LW-01",
    "rv32i_m/I/OR-01",
    "rv32i_m/I/ORI-01",
    "rv32i_m/I/SB-01",
    "rv32i_m/I/SH-01",
    "rv32i_m/I/SLL-01",
    "rv32i_m/I/SLLI-01",
    "rv32i_m/I/SLT-01",
    "rv32i_m/I/SLTI-01",
    "rv32i_m/I/SLTIU-01",
    "rv32i_m/I/SLTU-01",
    "rv32i_m/I/SRA-01",
    "rv32i_m/I/SRAI-01",
    "rv32i_m/I/SRL-01",
    "rv32i_m/I/SRLI-01",
    "rv32i_m/I/SUB-01",
    "rv32i_m/I/SW-01",
    "rv32i_m/I/XOR-01",
    "rv32i_m/I/XORI-01"   
  };

  string testsBP64[] = '{
    `IMPERASTEST,
    "rv64BP/simple",
    "rv64BP/mmm",
    "rv64BP/linpack_bench",
    "rv64BP/sieve",
    "rv64BP/qsort",
    "rv64BP/dhrystone"
  };

  string imperas32p[] = '{
    `MYIMPERASTEST,
    "rv32p/WALLY-MSTATUS",
    "rv32p/WALLY-MCAUSE",
    "rv32p/WALLY-SCAUSE",
    "rv32p/WALLY-MEPC",
    "rv32p/WALLY-SEPC",
    "rv32p/WALLY-MTVAL",
    "rv32p/WALLY-STVAL",
    "rv32p/WALLY-MARCHID",
    "rv32p/WALLY-MIMPID",
    "rv32p/WALLY-MHARTID",
    "rv32p/WALLY-MVENDORID",
    "rv32p/WALLY-MTVEC",
    "rv32p/WALLY-STVEC",
    "rv32p/WALLY-MIE",
    "rv32p/WALLY-MEDELEG",
    "rv32p/WALLY-IP",
    "rv32p/WALLY-CSR-PERMISSIONS-M",
    "rv32p/WALLY-CSR-PERMISSIONS-S"
  };

  string arch64priv[] = '{
    `RISCVARCHTEST,
    "rv64i_m/privilege/src/ebreak.S/ref/ref",
    "rv64i_m/privilege/src/ecall.S/ref/ref",
    "rv64i_m/privilege/src/misalign1-jalr-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign2-jalr-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-beq-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-bge-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-bgeu-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-blt-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-bltu-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-bne-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-jal-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-ld-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-lh-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-lhu-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-lw-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-lwu-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-sd-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-sh-01.S/ref/ref",
    "rv64i_m/privilege/src/misalign-sw-01.S/ref/ref"
    };

  string arch64m[] = '{
    `RISCVARCHTEST,
    "rv64i_m/M/src/div-01.S/ref/ref",
    "rv64i_m/M/src/divu-01.S/ref/ref",
    "rv64i_m/M/src/divuw-01.S/ref/ref",
    "rv64i_m/M/src/divw-01.S/ref/ref",
    "rv64i_m/M/src/mul-01.S/ref/ref",
    "rv64i_m/M/src/mulh-01.S/ref/ref",
    "rv64i_m/M/src/mulhsu-01.S/ref/ref",
    "rv64i_m/M/src/mulhu-01.S/ref/ref",
    "rv64i_m/M/src/mulw-01.S/ref/ref",
    "rv64i_m/M/src/rem-01.S/ref/ref",
    "rv64i_m/M/src/remu-01.S/ref/ref",
    "rv64i_m/M/src/remuw-01.S/ref/ref",
    "rv64i_m/M/src/remw-01.S/ref/ref"
   };

  string arch64c[] = '{
    `RISCVARCHTEST,
    "rv64i_m/C/src/cadd-01.S/ref/ref",
    "rv64i_m/C/src/caddi-01.S/ref/ref",
    "rv64i_m/C/src/caddi16sp-01.S/ref/ref",
    "rv64i_m/C/src/caddi4spn-01.S/ref/ref",
    "rv64i_m/C/src/caddiw-01.S/ref/ref",
    "rv64i_m/C/src/caddw-01.S/ref/ref",
    "rv64i_m/C/src/cand-01.S/ref/ref",
    "rv64i_m/C/src/candi-01.S/ref/ref",
    "rv64i_m/C/src/cbeqz-01.S/ref/ref",
    "rv64i_m/C/src/cbnez-01.S/ref/ref",
    "rv64i_m/C/src/cj-01.S/ref/ref",
    "rv64i_m/C/src/cjalr-01.S/ref/ref",
    "rv64i_m/C/src/cjr-01.S/ref/ref",
    "rv64i_m/C/src/cld-01.S/ref/ref",
    "rv64i_m/C/src/cldsp-01.S/ref/ref",
    "rv64i_m/C/src/cli-01.S/ref/ref",
    "rv64i_m/C/src/clui-01.S/ref/ref",
    "rv64i_m/C/src/clw-01.S/ref/ref",
    "rv64i_m/C/src/clwsp-01.S/ref/ref",
    "rv64i_m/C/src/cmv-01.S/ref/ref",
    "rv64i_m/C/src/cnop-01.S/ref/ref",
    "rv64i_m/C/src/cor-01.S/ref/ref",
    "rv64i_m/C/src/csd-01.S/ref/ref",
    "rv64i_m/C/src/csdsp-01.S/ref/ref",
    "rv64i_m/C/src/cslli-01.S/ref/ref",
    "rv64i_m/C/src/csrai-01.S/ref/ref",
    "rv64i_m/C/src/csrli-01.S/ref/ref",
    "rv64i_m/C/src/csub-01.S/ref/ref",
    "rv64i_m/C/src/csubw-01.S/ref/ref",
    "rv64i_m/C/src/csw-01.S/ref/ref",
    "rv64i_m/C/src/cswsp-01.S/ref/ref",
    "rv64i_m/C/src/cxor-01.S/ref/ref"
  };

  string arch64cpriv[] = '{
//    `RISCVARCHTEST,
    "rv64i_m/C/src/cebreak-01.S/ref/ref"
  };

  string arch64i[] = '{
    `RISCVARCHTEST,
    "rv64i_m/I/src/add-01.S/ref/ref",
    "rv64i_m/I/src/addi-01.S/ref/ref",
    "rv64i_m/I/src/addiw-01.S/ref/ref",
    "rv64i_m/I/src/addw-01.S/ref/ref",
    "rv64i_m/I/src/and-01.S/ref/ref",
    "rv64i_m/I/src/andi-01.S/ref/ref",
    "rv64i_m/I/src/auipc-01.S/ref/ref",
    "rv64i_m/I/src/beq-01.S/ref/ref",
    "rv64i_m/I/src/bge-01.S/ref/ref",
    "rv64i_m/I/src/bgeu-01.S/ref/ref",
    "rv64i_m/I/src/blt-01.S/ref/ref",
    "rv64i_m/I/src/bltu-01.S/ref/ref",
    "rv64i_m/I/src/bne-01.S/ref/ref",
    "rv64i_m/I/src/fence-01.S/ref/ref",
    "rv64i_m/I/src/jal-01.S/ref/ref",
    "rv64i_m/I/src/jalr-01.S/ref/ref",
    "rv64i_m/I/src/lb-align-01.S/ref/ref",
    "rv64i_m/I/src/lbu-align-01.S/ref/ref",
    "rv64i_m/I/src/ld-align-01.S/ref/ref",
    "rv64i_m/I/src/lh-align-01.S/ref/ref",
    "rv64i_m/I/src/lhu-align-01.S/ref/ref",
    "rv64i_m/I/src/lui-01.S/ref/ref",
    "rv64i_m/I/src/lw-align-01.S/ref/ref",
    "rv64i_m/I/src/lwu-align-01.S/ref/ref",
    "rv64i_m/I/src/or-01.S/ref/ref",
    "rv64i_m/I/src/ori-01.S/ref/ref",
    "rv64i_m/I/src/sb-align-01.S/ref/ref",
    "rv64i_m/I/src/sd-align-01.S/ref/ref",
    "rv64i_m/I/src/sh-align-01.S/ref/ref",
    "rv64i_m/I/src/sll-01.S/ref/ref",
    "rv64i_m/I/src/slli-01.S/ref/ref",
    "rv64i_m/I/src/slliw-01.S/ref/ref",
    "rv64i_m/I/src/sllw-01.S/ref/ref",
    "rv64i_m/I/src/slt-01.S/ref/ref",
    "rv64i_m/I/src/slti-01.S/ref/ref",
    "rv64i_m/I/src/sltiu-01.S/ref/ref",
    "rv64i_m/I/src/sltu-01.S/ref/ref",
    "rv64i_m/I/src/sra-01.S/ref/ref",
    "rv64i_m/I/src/srai-01.S/ref/ref",
    "rv64i_m/I/src/sraiw-01.S/ref/ref",
    "rv64i_m/I/src/sraw-01.S/ref/ref",
    "rv64i_m/I/src/srl-01.S/ref/ref",
    "rv64i_m/I/src/srli-01.S/ref/ref",
    "rv64i_m/I/src/srliw-01.S/ref/ref",
    "rv64i_m/I/src/srlw-01.S/ref/ref",
    "rv64i_m/I/src/sub-01.S/ref/ref",
    "rv64i_m/I/src/subw-01.S/ref/ref",
    "rv64i_m/I/src/sw-align-01.S/ref/ref",
    "rv64i_m/I/src/xor-01.S/ref/ref",
    "rv64i_m/I/src/xori-01.S/ref/ref"
  };

  string arch64d[] = '{
    `RISCVARCHTEST,
    "rv64i_m/D/src/d_fadd_b10-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b11-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b12-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b13-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fadd_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fclass_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.l_b25-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.l_b26-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.lu_b25-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.lu_b26-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.s_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.w_b25-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.w_b26-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.wu_b25-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.d.wu_b26-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.l.d_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.lu.d_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.s.d_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.w.d_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fcvt.wu.d_b29-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b1-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b20-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b2-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b21-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b3-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b4-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b5-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b6-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b7-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b8-01.S/ref/ref",
    // "rv64i_m/D/src/d_fdiv_b9-01.S/ref/ref",
    "rv64i_m/D/src/d_feq_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_feq_b19-01.S/ref/ref",
    "rv64i_m/D/src/d_fle_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fle_b19-01.S/ref/ref",
    "rv64i_m/D/src/d_flt_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_flt_b19-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b14-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b16-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b17-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b18-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b6-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fmadd_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fmax_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fmax_b19-01.S/ref/ref",
    "rv64i_m/D/src/d_fmin_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fmin_b19-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b14-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b16-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b17-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b18-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b6-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fmsub_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b6-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fmul_b9-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.d.x_b25-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.d.x_b26-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b22-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b23-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b24-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b27-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b28-01.S/ref/ref",
    "rv64i_m/D/src/d_fmv.x.d_b29-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b14-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b16-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b17-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b18-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b6-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmadd_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b14-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b16-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b17-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b18-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b6-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fnmsub_b8-01.S/ref/ref",
    "rv64i_m/D/src/d_fsgnj_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fsgnjn_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fsgnjx_b1-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b1-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b20-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b2-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b3-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b4-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b5-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b7-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b8-01.S/ref/ref",
    // "rv64i_m/D/src/d_fsqrt_b9-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b10-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b1-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b11-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b12-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b13-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b2-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b3-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b4-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b5-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b7-01.S/ref/ref",
    "rv64i_m/D/src/d_fsub_b8-01.S/ref/ref"
};

    string arch32priv[] = '{
    `RISCVARCHTEST,
    "rv32i_m/privilege/src/ebreak.S/ref/ref",
    "rv32i_m/privilege/src/ecall.S/ref/ref",
    "rv32i_m/privilege/src/misalign1-jalr-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign2-jalr-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-beq-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-bge-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-bgeu-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-blt-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-bltu-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-bne-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-jal-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-lh-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-lhu-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-lw-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-sh-01.S/ref/ref",
    "rv32i_m/privilege/src/misalign-sw-01.S/ref/ref"
    };

  string arch32m[] = '{
    `RISCVARCHTEST,
    "rv32i_m/M/src/div-01.S/ref/ref",
    "rv32i_m/M/src/divu-01.S/ref/ref",
    "rv32i_m/M/src/mul-01.S/ref/ref",
    "rv32i_m/M/src/mulh-01.S/ref/ref",
    "rv32i_m/M/src/mulhsu-01.S/ref/ref",
    "rv32i_m/M/src/mulhu-01.S/ref/ref",
    "rv32i_m/M/src/rem-01.S/ref/ref",
    "rv32i_m/M/src/remu-01.S/ref/ref"
   };

  string arch32f[] = '{
    `RISCVARCHTEST,
    "rv32i_m/F/src/fadd_b10-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b1-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b11-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b12-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b13-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b2-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b3-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b4-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b5-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b7-01.S/ref/ref",
    "rv32i_m/F/src/fadd_b8-01.S/ref/ref",
    "rv32i_m/F/src/fclass_b1-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.s.w_b25-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.s.w_b26-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.s.wu_b25-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.s.wu_b26-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b1-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b22-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b23-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b24-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b27-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b28-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.w.s_b29-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b1-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b22-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b23-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b24-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b27-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b28-01.S/ref/ref",
    "rv32i_m/F/src/fcvt.wu.s_b29-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b1-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b20-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b2-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b21-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b3-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b4-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b5-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b6-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b7-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b8-01.S/ref/ref",
    // "rv32i_m/F/src/fdiv_b9-01.S/ref/ref",
    "rv32i_m/F/src/feq_b1-01.S/ref/ref",
    "rv32i_m/F/src/feq_b19-01.S/ref/ref",
    "rv32i_m/F/src/fle_b1-01.S/ref/ref",
    "rv32i_m/F/src/fle_b19-01.S/ref/ref",
    "rv32i_m/F/src/flt_b1-01.S/ref/ref",
    "rv32i_m/F/src/flt_b19-01.S/ref/ref",
    "rv32i_m/F/src/flw-align-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b14-01.S/ref/ref",
    // "rv32i_m/F/src/fmadd_b15-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b16-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b17-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b18-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b2-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b3-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b4-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b5-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b6-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b7-01.S/ref/ref",
    "rv32i_m/F/src/fmadd_b8-01.S/ref/ref",
    "rv32i_m/F/src/fmax_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmax_b19-01.S/ref/ref",
    "rv32i_m/F/src/fmin_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmin_b19-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b14-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b15-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b16-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b17-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b18-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b2-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b3-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b4-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b5-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b6-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b7-01.S/ref/ref",
    "rv32i_m/F/src/fmsub_b8-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b2-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b3-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b4-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b5-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b6-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b7-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b8-01.S/ref/ref",
    "rv32i_m/F/src/fmul_b9-01.S/ref/ref",
    "rv32i_m/F/src/fmv.w.x_b25-01.S/ref/ref",
    "rv32i_m/F/src/fmv.w.x_b26-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b1-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b22-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b23-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b24-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b27-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b28-01.S/ref/ref",
    "rv32i_m/F/src/fmv.x.w_b29-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b1-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b14-01.S/ref/ref",
    // "rv32i_m/F/src/fnmadd_b15-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b16-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b17-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b18-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b2-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b3-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b4-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b5-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b6-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b7-01.S/ref/ref",
    "rv32i_m/F/src/fnmadd_b8-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b1-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b14-01.S/ref/ref",
    // "rv32i_m/F/src/fnmsub_b15-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b16-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b17-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b18-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b2-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b3-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b4-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b5-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b6-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b7-01.S/ref/ref",
    "rv32i_m/F/src/fnmsub_b8-01.S/ref/ref",
    "rv32i_m/F/src/fsgnj_b1-01.S/ref/ref",
    "rv32i_m/F/src/fsgnjn_b1-01.S/ref/ref",
    "rv32i_m/F/src/fsgnjx_b1-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b1-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b20-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b2-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b3-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b4-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b5-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b7-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b8-01.S/ref/ref",
    // "rv32i_m/F/src/fsqrt_b9-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b10-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b1-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b11-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b12-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b13-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b2-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b3-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b4-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b5-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b7-01.S/ref/ref",
    "rv32i_m/F/src/fsub_b8-01.S/ref/ref",
    "rv32i_m/F/src/fsw-align-01.S/ref/ref"
    };


  string arch32c[] = '{
    `RISCVARCHTEST,
    "rv32i_m/C/src/cadd-01.S/ref/ref",
  "rv32i_m/C/src/caddi-01.S/ref/ref",
  "rv32i_m/C/src/caddi16sp-01.S/ref/ref",
  "rv32i_m/C/src/caddi4spn-01.S/ref/ref",
  "rv32i_m/C/src/cand-01.S/ref/ref",
  "rv32i_m/C/src/candi-01.S/ref/ref",
  "rv32i_m/C/src/cbeqz-01.S/ref/ref",
  "rv32i_m/C/src/cbnez-01.S/ref/ref",
  "rv32i_m/C/src/cj-01.S/ref/ref",
  "rv32i_m/C/src/cjal-01.S/ref/ref",
  "rv32i_m/C/src/cjalr-01.S/ref/ref",
  "rv32i_m/C/src/cjr-01.S/ref/ref",
  "rv32i_m/C/src/cli-01.S/ref/ref",
  "rv32i_m/C/src/clui-01.S/ref/ref",
  "rv32i_m/C/src/clw-01.S/ref/ref",
  "rv32i_m/C/src/clwsp-01.S/ref/ref",
  "rv32i_m/C/src/cmv-01.S/ref/ref",
  "rv32i_m/C/src/cnop-01.S/ref/ref",
  "rv32i_m/C/src/cor-01.S/ref/ref",
  "rv32i_m/C/src/cslli-01.S/ref/ref",
  "rv32i_m/C/src/csrai-01.S/ref/ref",
  "rv32i_m/C/src/csrli-01.S/ref/ref",
  "rv32i_m/C/src/csub-01.S/ref/ref",
  "rv32i_m/C/src/csw-01.S/ref/ref",
  "rv32i_m/C/src/cswsp-01.S/ref/ref",
  "rv32i_m/C/src/cxor-01.S/ref/ref"
  };

  string arch32cpriv[] = '{
  //  `RISCVARCHTEST,
  "rv32i_m/C/src/cebreak-01.S/ref/ref"
  };      


  string arch32i[] = '{
    `RISCVARCHTEST,
    "rv32i_m/I/src/add-01.S/ref/ref",
    "rv32i_m/I/src/addi-01.S/ref/ref",
    "rv32i_m/I/src/and-01.S/ref/ref",
    "rv32i_m/I/src/andi-01.S/ref/ref",
    "rv32i_m/I/src/auipc-01.S/ref/ref",
    "rv32i_m/I/src/beq-01.S/ref/ref",
    "rv32i_m/I/src/bge-01.S/ref/ref",
    "rv32i_m/I/src/bgeu-01.S/ref/ref",
    "rv32i_m/I/src/blt-01.S/ref/ref",
    "rv32i_m/I/src/bltu-01.S/ref/ref",
    "rv32i_m/I/src/bne-01.S/ref/ref",
    "rv32i_m/I/src/fence-01.S/ref/ref",
    "rv32i_m/I/src/jal-01.S/ref/ref",
    "rv32i_m/I/src/jalr-01.S/ref/ref",
    "rv32i_m/I/src/lb-align-01.S/ref/ref",
    "rv32i_m/I/src/lbu-align-01.S/ref/ref",
    "rv32i_m/I/src/lh-align-01.S/ref/ref",
    "rv32i_m/I/src/lhu-align-01.S/ref/ref",
    "rv32i_m/I/src/lui-01.S/ref/ref",
    "rv32i_m/I/src/lw-align-01.S/ref/ref",
    "rv32i_m/I/src/or-01.S/ref/ref",
    "rv32i_m/I/src/ori-01.S/ref/ref",
    "rv32i_m/I/src/sb-align-01.S/ref/ref",
    "rv32i_m/I/src/sh-align-01.S/ref/ref",
    "rv32i_m/I/src/sll-01.S/ref/ref",
    "rv32i_m/I/src/slli-01.S/ref/ref",
    "rv32i_m/I/src/slt-01.S/ref/ref",
    "rv32i_m/I/src/slti-01.S/ref/ref",
    "rv32i_m/I/src/sltiu-01.S/ref/ref",
    "rv32i_m/I/src/sltu-01.S/ref/ref",
    "rv32i_m/I/src/sra-01.S/ref/ref",
    "rv32i_m/I/src/srai-01.S/ref/ref",
    "rv32i_m/I/src/srl-01.S/ref/ref",
    "rv32i_m/I/src/srli-01.S/ref/ref",
    "rv32i_m/I/src/sub-01.S/ref/ref",
    "rv32i_m/I/src/sw-align-01.S/ref/ref",
    "rv32i_m/I/src/xor-01.S/ref/ref",
    "rv32i_m/I/src/xori-01.S/ref/ref"
  };

 string wally64i[] = '{
    `WALLYTEST,
    "rv64i_m/I/WALLY-ADD",
    "rv64i_m/I/WALLY-SLT",
    "rv64i_m/I/WALLY-SLTU",
    "rv64i_m/I/WALLY-SUB",
    "rv64i_m/I/WALLY-XOR"
 };

 string wally64priv[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-status-tw-01",
    "rv64i_m/privilege/WALLY-csr-permission-s-01",
    "rv64i_m/privilege/WALLY-csr-permission-u-01",
    "rv64i_m/privilege/WALLY-minfo-01",
    "rv64i_m/privilege/WALLY-misa-01",
    "rv64i_m/privilege/WALLY-mmu-sv39",
    "rv64i_m/privilege/WALLY-mmu-sv48",
    "rv64i_m/privilege/WALLY-pma",
    "rv64i_m/privilege/WALLY-pmp",
    "rv64i_m/privilege/WALLY-trap-01",
    "rv64i_m/privilege/WALLY-trap-s-01",
    "rv64i_m/privilege/WALLY-trap-u-01",
    "rv64i_m/privilege/WALLY-mie-01",
    "rv64i_m/privilege/WALLY-sie-01",
    "rv64i_m/privilege/WALLY-mtvec-01",
    "rv64i_m/privilege/WALLY-stvec-01",
    "rv64i_m/privilege/WALLY-status-mie-01",
    "rv64i_m/privilege/WALLY-status-sie-01",
    "rv64i_m/privilege/WALLY-trap-sret-01",
    "rv64i_m/privilege/WALLY-status-tw-01",
    "rv64i_m/privilege/WALLY-wfi-01"
 };

 string wally64periph[] = '{
    `WALLYTEST,
    "rv64i_m/privilege/WALLY-periph"
 };

 string wally32e[] = '{
    `WALLYTEST,
    "rv32i_m/I/E-add-01",
    "rv32i_m/I/E-addi-01",
    "rv32i_m/I/E-and-01",
    "rv32i_m/I/E-andi-01",
    "rv32i_m/I/E-auipc-01",
    "rv32i_m/I/E-bge-01",
    "rv32i_m/I/E-bgeu-01",
    "rv32i_m/I/E-blt-01",
    "rv32i_m/I/E-bltu-01",
    "rv32i_m/I/E-bne-01",
    "rv32i_m/I/E-jal-01",
    "rv32i_m/I/E-jalr-01",
    "rv32i_m/I/E-lb-align-01",
    "rv32i_m/I/E-lbu-align-01",
    "rv32i_m/I/E-lh-align-01",
    "rv32i_m/I/E-lhu-align-01",
    "rv32i_m/I/E-lui-01",
    "rv32i_m/I/E-lw-align-01",
    "rv32i_m/I/E-or-01",
    "rv32i_m/I/E-ori-01",
    "rv32i_m/I/E-sb-align-01",
    "rv32i_m/I/E-sh-align-01",
    "rv32i_m/I/E-sll-01",
    "rv32i_m/I/E-slli-01",
    "rv32i_m/I/E-slt-01",
    "rv32i_m/I/E-slti-01",
    "rv32i_m/I/E-sltiu-01",
    "rv32i_m/I/E-sltu-01",
    "rv32i_m/I/E-sra-01",
    "rv32i_m/I/E-srai-01",
    "rv32i_m/I/E-srl-01",
    "rv32i_m/I/E-srli-01",
    "rv32i_m/I/E-sub-01",
    "rv32i_m/I/E-sw-align-01",
    "rv32i_m/I/E-xor-01",
    "rv32i_m/I/E-xori-01"
 };

string wally32i[] = '{
    `WALLYTEST,
    "rv32i_m/I/WALLY-ADD",
    "rv32i_m/I/WALLY-SLT",
    "rv32i_m/I/WALLY-SLTU",
    "rv32i_m/I/WALLY-SUB",
    "rv32i_m/I/WALLY-XOR"
 };

 string wally32priv[] = '{
    `WALLYTEST,
    "rv32i_m/privilege/WALLY-csr-permission-s-01",
    "rv32i_m/privilege/WALLY-csr-permission-u-01",
    "rv32i_m/privilege/WALLY-minfo-01",
    "rv32i_m/privilege/WALLY-misa-01",
    "rv32i_m/privilege/WALLY-mmu-sv32",
    "rv32i_m/privilege/WALLY-pma",
    "rv32i_m/privilege/WALLY-pmp",
    "rv32i_m/privilege/WALLY-trap-01",
    "rv32i_m/privilege/WALLY-trap-s-01",
    "rv32i_m/privilege/WALLY-trap-u-01",
    "rv32i_m/privilege/WALLY-mie-01",
    "rv32i_m/privilege/WALLY-sie-01",
    "rv32i_m/privilege/WALLY-mtvec-01",
    "rv32i_m/privilege/WALLY-stvec-01",
    "rv32i_m/privilege/WALLY-status-mie-01",
    "rv32i_m/privilege/WALLY-status-sie-01",
    "rv32i_m/privilege/WALLY-trap-sret-01",
    "rv32i_m/privilege/WALLY-status-tw-01", 
    "rv32i_m/privilege/WALLY-wfi-01"
 };

 string wally32periph[] = '{
    `WALLYTEST
 };


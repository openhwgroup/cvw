test_fencei_cg = new(); test_fencei_cg.set_inst_name("obj_fencei");

//    test_fencei_cg = new(); 
//test_fencei_cg.set_inst_name("obj_fencei");

../../../config/rv32gc/coverage.svh
// James Kaden Cassidy
// kacassidy@hmc.edu
// 1/5/2026

`ifndef PARAMETERS
`define PARAMETERS

    `define XLEN 32

    //`define DEBUG

`endif
